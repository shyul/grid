// frontier.v

// Generated using ACDS version 11.1sp2 259 at 2012.07.20.15:59:36

`timescale 1 ps / 1 ps
module frontier (
		input  wire        a20_f0_oe,      //    a20.f0_oe
		input  wire        a20_f1_oe,      //       .f1_oe
		input  wire        a20_f2_oe,      //       .f2_oe
		input  wire        a20_f3_oe,      //       .f3_oe
		input  wire        a20_f4_oe,      //       .f4_oe
		input  wire        a20_f5_oe,      //       .f5_oe
		input  wire        a20_f6_oe,      //       .f6_oe
		input  wire        a20_f7_oe,      //       .f7_oe
		input  wire        a20_f0_out,     //       .f0_out
		input  wire        a20_f1_out,     //       .f1_out
		input  wire        a20_f2_out,     //       .f2_out
		input  wire        a20_f3_out,     //       .f3_out
		input  wire        a20_f4_out,     //       .f4_out
		input  wire        a20_f5_out,     //       .f5_out
		input  wire        a20_f6_out,     //       .f6_out
		input  wire        a20_f7_out,     //       .f7_out
		output wire        a20_f_in,       //       .f_in
		inout  wire        a20_GPIO,       //       .GPIO
		input  wire        b19_f0_oe,      //    b19.f0_oe
		input  wire        b19_f1_oe,      //       .f1_oe
		input  wire        b19_f2_oe,      //       .f2_oe
		input  wire        b19_f3_oe,      //       .f3_oe
		input  wire        b19_f4_oe,      //       .f4_oe
		input  wire        b19_f5_oe,      //       .f5_oe
		input  wire        b19_f6_oe,      //       .f6_oe
		input  wire        b19_f7_oe,      //       .f7_oe
		input  wire        b19_f0_out,     //       .f0_out
		input  wire        b19_f1_out,     //       .f1_out
		input  wire        b19_f2_out,     //       .f2_out
		input  wire        b19_f3_out,     //       .f3_out
		input  wire        b19_f4_out,     //       .f4_out
		input  wire        b19_f5_out,     //       .f5_out
		input  wire        b19_f6_out,     //       .f6_out
		input  wire        b19_f7_out,     //       .f7_out
		output wire        b19_f_in,       //       .f_in
		inout  wire        b19_GPIO,       //       .GPIO
		input  wire        a16_f0_oe,      //    a16.f0_oe
		input  wire        a16_f1_oe,      //       .f1_oe
		input  wire        a16_f2_oe,      //       .f2_oe
		input  wire        a16_f3_oe,      //       .f3_oe
		input  wire        a16_f4_oe,      //       .f4_oe
		input  wire        a16_f5_oe,      //       .f5_oe
		input  wire        a16_f6_oe,      //       .f6_oe
		input  wire        a16_f7_oe,      //       .f7_oe
		input  wire        a16_f0_out,     //       .f0_out
		input  wire        a16_f1_out,     //       .f1_out
		input  wire        a16_f2_out,     //       .f2_out
		input  wire        a16_f3_out,     //       .f3_out
		input  wire        a16_f4_out,     //       .f4_out
		input  wire        a16_f5_out,     //       .f5_out
		input  wire        a16_f6_out,     //       .f6_out
		input  wire        a16_f7_out,     //       .f7_out
		output wire        a16_f_in,       //       .f_in
		inout  wire        a16_GPIO,       //       .GPIO
		input  wire        a17_f0_oe,      //    a17.f0_oe
		input  wire        a17_f1_oe,      //       .f1_oe
		input  wire        a17_f2_oe,      //       .f2_oe
		input  wire        a17_f3_oe,      //       .f3_oe
		input  wire        a17_f4_oe,      //       .f4_oe
		input  wire        a17_f5_oe,      //       .f5_oe
		input  wire        a17_f6_oe,      //       .f6_oe
		input  wire        a17_f7_oe,      //       .f7_oe
		input  wire        a17_f0_out,     //       .f0_out
		input  wire        a17_f1_out,     //       .f1_out
		input  wire        a17_f2_out,     //       .f2_out
		input  wire        a17_f3_out,     //       .f3_out
		input  wire        a17_f4_out,     //       .f4_out
		input  wire        a17_f5_out,     //       .f5_out
		input  wire        a17_f6_out,     //       .f6_out
		input  wire        a17_f7_out,     //       .f7_out
		output wire        a17_f_in,       //       .f_in
		inout  wire        a17_GPIO,       //       .GPIO
		input  wire        b17_f0_oe,      //    b17.f0_oe
		input  wire        b17_f1_oe,      //       .f1_oe
		input  wire        b17_f2_oe,      //       .f2_oe
		input  wire        b17_f3_oe,      //       .f3_oe
		input  wire        b17_f4_oe,      //       .f4_oe
		input  wire        b17_f5_oe,      //       .f5_oe
		input  wire        b17_f6_oe,      //       .f6_oe
		input  wire        b17_f7_oe,      //       .f7_oe
		input  wire        b17_f0_out,     //       .f0_out
		input  wire        b17_f1_out,     //       .f1_out
		input  wire        b17_f2_out,     //       .f2_out
		input  wire        b17_f3_out,     //       .f3_out
		input  wire        b17_f4_out,     //       .f4_out
		input  wire        b17_f5_out,     //       .f5_out
		input  wire        b17_f6_out,     //       .f6_out
		input  wire        b17_f7_out,     //       .f7_out
		output wire        b17_f_in,       //       .f_in
		inout  wire        b17_GPIO,       //       .GPIO
		input  wire        a14_f0_oe,      //    a14.f0_oe
		input  wire        a14_f1_oe,      //       .f1_oe
		input  wire        a14_f2_oe,      //       .f2_oe
		input  wire        a14_f3_oe,      //       .f3_oe
		input  wire        a14_f4_oe,      //       .f4_oe
		input  wire        a14_f5_oe,      //       .f5_oe
		input  wire        a14_f6_oe,      //       .f6_oe
		input  wire        a14_f7_oe,      //       .f7_oe
		input  wire        a14_f0_out,     //       .f0_out
		input  wire        a14_f1_out,     //       .f1_out
		input  wire        a14_f2_out,     //       .f2_out
		input  wire        a14_f3_out,     //       .f3_out
		input  wire        a14_f4_out,     //       .f4_out
		input  wire        a14_f5_out,     //       .f5_out
		input  wire        a14_f6_out,     //       .f6_out
		input  wire        a14_f7_out,     //       .f7_out
		output wire        a14_f_in,       //       .f_in
		inout  wire        a14_GPIO,       //       .GPIO
		input  wire        b18_f0_oe,      //    b18.f0_oe
		input  wire        b18_f1_oe,      //       .f1_oe
		input  wire        b18_f2_oe,      //       .f2_oe
		input  wire        b18_f3_oe,      //       .f3_oe
		input  wire        b18_f4_oe,      //       .f4_oe
		input  wire        b18_f5_oe,      //       .f5_oe
		input  wire        b18_f6_oe,      //       .f6_oe
		input  wire        b18_f7_oe,      //       .f7_oe
		input  wire        b18_f0_out,     //       .f0_out
		input  wire        b18_f1_out,     //       .f1_out
		input  wire        b18_f2_out,     //       .f2_out
		input  wire        b18_f3_out,     //       .f3_out
		input  wire        b18_f4_out,     //       .f4_out
		input  wire        b18_f5_out,     //       .f5_out
		input  wire        b18_f6_out,     //       .f6_out
		input  wire        b18_f7_out,     //       .f7_out
		output wire        b18_f_in,       //       .f_in
		inout  wire        b18_GPIO,       //       .GPIO
		input  wire        a15_f0_oe,      //    a15.f0_oe
		input  wire        a15_f1_oe,      //       .f1_oe
		input  wire        a15_f2_oe,      //       .f2_oe
		input  wire        a15_f3_oe,      //       .f3_oe
		input  wire        a15_f4_oe,      //       .f4_oe
		input  wire        a15_f5_oe,      //       .f5_oe
		input  wire        a15_f6_oe,      //       .f6_oe
		input  wire        a15_f7_oe,      //       .f7_oe
		input  wire        a15_f0_out,     //       .f0_out
		input  wire        a15_f1_out,     //       .f1_out
		input  wire        a15_f2_out,     //       .f2_out
		input  wire        a15_f3_out,     //       .f3_out
		input  wire        a15_f4_out,     //       .f4_out
		input  wire        a15_f5_out,     //       .f5_out
		input  wire        a15_f6_out,     //       .f6_out
		input  wire        a15_f7_out,     //       .f7_out
		output wire        a15_f_in,       //       .f_in
		inout  wire        a15_GPIO,       //       .GPIO
		input  wire        a12_f0_oe,      //    a12.f0_oe
		input  wire        a12_f1_oe,      //       .f1_oe
		input  wire        a12_f2_oe,      //       .f2_oe
		input  wire        a12_f3_oe,      //       .f3_oe
		input  wire        a12_f4_oe,      //       .f4_oe
		input  wire        a12_f5_oe,      //       .f5_oe
		input  wire        a12_f6_oe,      //       .f6_oe
		input  wire        a12_f7_oe,      //       .f7_oe
		input  wire        a12_f0_out,     //       .f0_out
		input  wire        a12_f1_out,     //       .f1_out
		input  wire        a12_f2_out,     //       .f2_out
		input  wire        a12_f3_out,     //       .f3_out
		input  wire        a12_f4_out,     //       .f4_out
		input  wire        a12_f5_out,     //       .f5_out
		input  wire        a12_f6_out,     //       .f6_out
		input  wire        a12_f7_out,     //       .f7_out
		output wire        a12_f_in,       //       .f_in
		inout  wire        a12_GPIO,       //       .GPIO
		input  wire        a13_f0_oe,      //    a13.f0_oe
		input  wire        a13_f1_oe,      //       .f1_oe
		input  wire        a13_f2_oe,      //       .f2_oe
		input  wire        a13_f3_oe,      //       .f3_oe
		input  wire        a13_f4_oe,      //       .f4_oe
		input  wire        a13_f5_oe,      //       .f5_oe
		input  wire        a13_f6_oe,      //       .f6_oe
		input  wire        a13_f7_oe,      //       .f7_oe
		input  wire        a13_f0_out,     //       .f0_out
		input  wire        a13_f1_out,     //       .f1_out
		input  wire        a13_f2_out,     //       .f2_out
		input  wire        a13_f3_out,     //       .f3_out
		input  wire        a13_f4_out,     //       .f4_out
		input  wire        a13_f5_out,     //       .f5_out
		input  wire        a13_f6_out,     //       .f6_out
		input  wire        a13_f7_out,     //       .f7_out
		output wire        a13_f_in,       //       .f_in
		inout  wire        a13_GPIO,       //       .GPIO
		input  wire        a10_f0_oe,      //    a10.f0_oe
		input  wire        a10_f1_oe,      //       .f1_oe
		input  wire        a10_f2_oe,      //       .f2_oe
		input  wire        a10_f3_oe,      //       .f3_oe
		input  wire        a10_f4_oe,      //       .f4_oe
		input  wire        a10_f5_oe,      //       .f5_oe
		input  wire        a10_f6_oe,      //       .f6_oe
		input  wire        a10_f7_oe,      //       .f7_oe
		input  wire        a10_f0_out,     //       .f0_out
		input  wire        a10_f1_out,     //       .f1_out
		input  wire        a10_f2_out,     //       .f2_out
		input  wire        a10_f3_out,     //       .f3_out
		input  wire        a10_f4_out,     //       .f4_out
		input  wire        a10_f5_out,     //       .f5_out
		input  wire        a10_f6_out,     //       .f6_out
		input  wire        a10_f7_out,     //       .f7_out
		output wire        a10_f_in,       //       .f_in
		inout  wire        a10_GPIO,       //       .GPIO
		input  wire        a11_f0_oe,      //    a11.f0_oe
		input  wire        a11_f1_oe,      //       .f1_oe
		input  wire        a11_f2_oe,      //       .f2_oe
		input  wire        a11_f3_oe,      //       .f3_oe
		input  wire        a11_f4_oe,      //       .f4_oe
		input  wire        a11_f5_oe,      //       .f5_oe
		input  wire        a11_f6_oe,      //       .f6_oe
		input  wire        a11_f7_oe,      //       .f7_oe
		input  wire        a11_f0_out,     //       .f0_out
		input  wire        a11_f1_out,     //       .f1_out
		input  wire        a11_f2_out,     //       .f2_out
		input  wire        a11_f3_out,     //       .f3_out
		input  wire        a11_f4_out,     //       .f4_out
		input  wire        a11_f5_out,     //       .f5_out
		input  wire        a11_f6_out,     //       .f6_out
		input  wire        a11_f7_out,     //       .f7_out
		output wire        a11_f_in,       //       .f_in
		inout  wire        a11_GPIO,       //       .GPIO
		input  wire        b11_f0_oe,      //    b11.f0_oe
		input  wire        b11_f1_oe,      //       .f1_oe
		input  wire        b11_f2_oe,      //       .f2_oe
		input  wire        b11_f3_oe,      //       .f3_oe
		input  wire        b11_f4_oe,      //       .f4_oe
		input  wire        b11_f5_oe,      //       .f5_oe
		input  wire        b11_f6_oe,      //       .f6_oe
		input  wire        b11_f7_oe,      //       .f7_oe
		input  wire        b11_f0_out,     //       .f0_out
		input  wire        b11_f1_out,     //       .f1_out
		input  wire        b11_f2_out,     //       .f2_out
		input  wire        b11_f3_out,     //       .f3_out
		input  wire        b11_f4_out,     //       .f4_out
		input  wire        b11_f5_out,     //       .f5_out
		input  wire        b11_f6_out,     //       .f6_out
		input  wire        b11_f7_out,     //       .f7_out
		output wire        b11_f_in,       //       .f_in
		inout  wire        b11_GPIO,       //       .GPIO
		input  wire        b12_f0_oe,      //    b12.f0_oe
		input  wire        b12_f1_oe,      //       .f1_oe
		input  wire        b12_f2_oe,      //       .f2_oe
		input  wire        b12_f3_oe,      //       .f3_oe
		input  wire        b12_f4_oe,      //       .f4_oe
		input  wire        b12_f5_oe,      //       .f5_oe
		input  wire        b12_f6_oe,      //       .f6_oe
		input  wire        b12_f7_oe,      //       .f7_oe
		input  wire        b12_f0_out,     //       .f0_out
		input  wire        b12_f1_out,     //       .f1_out
		input  wire        b12_f2_out,     //       .f2_out
		input  wire        b12_f3_out,     //       .f3_out
		input  wire        b12_f4_out,     //       .f4_out
		input  wire        b12_f5_out,     //       .f5_out
		input  wire        b12_f6_out,     //       .f6_out
		input  wire        b12_f7_out,     //       .f7_out
		output wire        b12_f_in,       //       .f_in
		inout  wire        b12_GPIO,       //       .GPIO
		input  wire        b10_f0_oe,      //    b10.f0_oe
		input  wire        b10_f1_oe,      //       .f1_oe
		input  wire        b10_f2_oe,      //       .f2_oe
		input  wire        b10_f3_oe,      //       .f3_oe
		input  wire        b10_f4_oe,      //       .f4_oe
		input  wire        b10_f5_oe,      //       .f5_oe
		input  wire        b10_f6_oe,      //       .f6_oe
		input  wire        b10_f7_oe,      //       .f7_oe
		input  wire        b10_f0_out,     //       .f0_out
		input  wire        b10_f1_out,     //       .f1_out
		input  wire        b10_f2_out,     //       .f2_out
		input  wire        b10_f3_out,     //       .f3_out
		input  wire        b10_f4_out,     //       .f4_out
		input  wire        b10_f5_out,     //       .f5_out
		input  wire        b10_f6_out,     //       .f6_out
		input  wire        b10_f7_out,     //       .f7_out
		output wire        b10_f_in,       //       .f_in
		inout  wire        b10_GPIO,       //       .GPIO
		input  wire        b15_f0_oe,      //    b15.f0_oe
		input  wire        b15_f1_oe,      //       .f1_oe
		input  wire        b15_f2_oe,      //       .f2_oe
		input  wire        b15_f3_oe,      //       .f3_oe
		input  wire        b15_f4_oe,      //       .f4_oe
		input  wire        b15_f5_oe,      //       .f5_oe
		input  wire        b15_f6_oe,      //       .f6_oe
		input  wire        b15_f7_oe,      //       .f7_oe
		input  wire        b15_f0_out,     //       .f0_out
		input  wire        b15_f1_out,     //       .f1_out
		input  wire        b15_f2_out,     //       .f2_out
		input  wire        b15_f3_out,     //       .f3_out
		input  wire        b15_f4_out,     //       .f4_out
		input  wire        b15_f5_out,     //       .f5_out
		input  wire        b15_f6_out,     //       .f6_out
		input  wire        b15_f7_out,     //       .f7_out
		output wire        b15_f_in,       //       .f_in
		inout  wire        b15_GPIO,       //       .GPIO
		input  wire        b16_f0_oe,      //    b16.f0_oe
		input  wire        b16_f1_oe,      //       .f1_oe
		input  wire        b16_f2_oe,      //       .f2_oe
		input  wire        b16_f3_oe,      //       .f3_oe
		input  wire        b16_f4_oe,      //       .f4_oe
		input  wire        b16_f5_oe,      //       .f5_oe
		input  wire        b16_f6_oe,      //       .f6_oe
		input  wire        b16_f7_oe,      //       .f7_oe
		input  wire        b16_f0_out,     //       .f0_out
		input  wire        b16_f1_out,     //       .f1_out
		input  wire        b16_f2_out,     //       .f2_out
		input  wire        b16_f3_out,     //       .f3_out
		input  wire        b16_f4_out,     //       .f4_out
		input  wire        b16_f5_out,     //       .f5_out
		input  wire        b16_f6_out,     //       .f6_out
		input  wire        b16_f7_out,     //       .f7_out
		output wire        b16_f_in,       //       .f_in
		inout  wire        b16_GPIO,       //       .GPIO
		input  wire        b13_f0_oe,      //    b13.f0_oe
		input  wire        b13_f1_oe,      //       .f1_oe
		input  wire        b13_f2_oe,      //       .f2_oe
		input  wire        b13_f3_oe,      //       .f3_oe
		input  wire        b13_f4_oe,      //       .f4_oe
		input  wire        b13_f5_oe,      //       .f5_oe
		input  wire        b13_f6_oe,      //       .f6_oe
		input  wire        b13_f7_oe,      //       .f7_oe
		input  wire        b13_f0_out,     //       .f0_out
		input  wire        b13_f1_out,     //       .f1_out
		input  wire        b13_f2_out,     //       .f2_out
		input  wire        b13_f3_out,     //       .f3_out
		input  wire        b13_f4_out,     //       .f4_out
		input  wire        b13_f5_out,     //       .f5_out
		input  wire        b13_f6_out,     //       .f6_out
		input  wire        b13_f7_out,     //       .f7_out
		output wire        b13_f_in,       //       .f_in
		inout  wire        b13_GPIO,       //       .GPIO
		input  wire        a18_f0_oe,      //    a18.f0_oe
		input  wire        a18_f1_oe,      //       .f1_oe
		input  wire        a18_f2_oe,      //       .f2_oe
		input  wire        a18_f3_oe,      //       .f3_oe
		input  wire        a18_f4_oe,      //       .f4_oe
		input  wire        a18_f5_oe,      //       .f5_oe
		input  wire        a18_f6_oe,      //       .f6_oe
		input  wire        a18_f7_oe,      //       .f7_oe
		input  wire        a18_f0_out,     //       .f0_out
		input  wire        a18_f1_out,     //       .f1_out
		input  wire        a18_f2_out,     //       .f2_out
		input  wire        a18_f3_out,     //       .f3_out
		input  wire        a18_f4_out,     //       .f4_out
		input  wire        a18_f5_out,     //       .f5_out
		input  wire        a18_f6_out,     //       .f6_out
		input  wire        a18_f7_out,     //       .f7_out
		output wire        a18_f_in,       //       .f_in
		inout  wire        a18_GPIO,       //       .GPIO
		input  wire        b14_f0_oe,      //    b14.f0_oe
		input  wire        b14_f1_oe,      //       .f1_oe
		input  wire        b14_f2_oe,      //       .f2_oe
		input  wire        b14_f3_oe,      //       .f3_oe
		input  wire        b14_f4_oe,      //       .f4_oe
		input  wire        b14_f5_oe,      //       .f5_oe
		input  wire        b14_f6_oe,      //       .f6_oe
		input  wire        b14_f7_oe,      //       .f7_oe
		input  wire        b14_f0_out,     //       .f0_out
		input  wire        b14_f1_out,     //       .f1_out
		input  wire        b14_f2_out,     //       .f2_out
		input  wire        b14_f3_out,     //       .f3_out
		input  wire        b14_f4_out,     //       .f4_out
		input  wire        b14_f5_out,     //       .f5_out
		input  wire        b14_f6_out,     //       .f6_out
		input  wire        b14_f7_out,     //       .f7_out
		output wire        b14_f_in,       //       .f_in
		inout  wire        b14_GPIO,       //       .GPIO
		input  wire        a19_f0_oe,      //    a19.f0_oe
		input  wire        a19_f1_oe,      //       .f1_oe
		input  wire        a19_f2_oe,      //       .f2_oe
		input  wire        a19_f3_oe,      //       .f3_oe
		input  wire        a19_f4_oe,      //       .f4_oe
		input  wire        a19_f5_oe,      //       .f5_oe
		input  wire        a19_f6_oe,      //       .f6_oe
		input  wire        a19_f7_oe,      //       .f7_oe
		input  wire        a19_f0_out,     //       .f0_out
		input  wire        a19_f1_out,     //       .f1_out
		input  wire        a19_f2_out,     //       .f2_out
		input  wire        a19_f3_out,     //       .f3_out
		input  wire        a19_f4_out,     //       .f4_out
		input  wire        a19_f5_out,     //       .f5_out
		input  wire        a19_f6_out,     //       .f6_out
		input  wire        a19_f7_out,     //       .f7_out
		output wire        a19_f_in,       //       .f_in
		inout  wire        a19_GPIO,       //       .GPIO
		input  wire        m1_RSTN,        //     m1.RSTN
		input  wire        m1_CLK,         //       .CLK
		input  wire [21:0] m1_ADDR,        //       .ADDR
		inout  wire [31:0] m1_DATA,        //       .DATA
		input  wire [3:0]  m1_CSN,         //       .CSN
		input  wire [3:0]  m1_BEN,         //       .BEN
		input  wire        m1_RDN,         //       .RDN
		input  wire        m1_WRN,         //       .WRN
		output wire        m1_WAITN,       //       .WAITN
		output wire [9:0]  m1_EINT,        //       .EINT
		input  wire        a25_f0_oe,      //    a25.f0_oe
		input  wire        a25_f1_oe,      //       .f1_oe
		input  wire        a25_f2_oe,      //       .f2_oe
		input  wire        a25_f3_oe,      //       .f3_oe
		input  wire        a25_f4_oe,      //       .f4_oe
		input  wire        a25_f5_oe,      //       .f5_oe
		input  wire        a25_f6_oe,      //       .f6_oe
		input  wire        a25_f7_oe,      //       .f7_oe
		input  wire        a25_f0_out,     //       .f0_out
		input  wire        a25_f1_out,     //       .f1_out
		input  wire        a25_f2_out,     //       .f2_out
		input  wire        a25_f3_out,     //       .f3_out
		input  wire        a25_f4_out,     //       .f4_out
		input  wire        a25_f5_out,     //       .f5_out
		input  wire        a25_f6_out,     //       .f6_out
		input  wire        a25_f7_out,     //       .f7_out
		output wire        a25_f_in,       //       .f_in
		inout  wire        a25_GPIO,       //       .GPIO
		output wire        led_f3_R,       // led_f3.R
		output wire        led_f3_G,       //       .G
		output wire        led_f3_B,       //       .B
		output wire        led_f2_R,       // led_f2.R
		output wire        led_f2_G,       //       .G
		output wire        led_f2_B,       //       .B
		input  wire        a21_f0_oe,      //    a21.f0_oe
		input  wire        a21_f1_oe,      //       .f1_oe
		input  wire        a21_f2_oe,      //       .f2_oe
		input  wire        a21_f3_oe,      //       .f3_oe
		input  wire        a21_f4_oe,      //       .f4_oe
		input  wire        a21_f5_oe,      //       .f5_oe
		input  wire        a21_f6_oe,      //       .f6_oe
		input  wire        a21_f7_oe,      //       .f7_oe
		input  wire        a21_f0_out,     //       .f0_out
		input  wire        a21_f1_out,     //       .f1_out
		input  wire        a21_f2_out,     //       .f2_out
		input  wire        a21_f3_out,     //       .f3_out
		input  wire        a21_f4_out,     //       .f4_out
		input  wire        a21_f5_out,     //       .f5_out
		input  wire        a21_f6_out,     //       .f6_out
		input  wire        a21_f7_out,     //       .f7_out
		output wire        a21_f_in,       //       .f_in
		inout  wire        a21_GPIO,       //       .GPIO
		input  wire        a22_f0_oe,      //    a22.f0_oe
		input  wire        a22_f1_oe,      //       .f1_oe
		input  wire        a22_f2_oe,      //       .f2_oe
		input  wire        a22_f3_oe,      //       .f3_oe
		input  wire        a22_f4_oe,      //       .f4_oe
		input  wire        a22_f5_oe,      //       .f5_oe
		input  wire        a22_f6_oe,      //       .f6_oe
		input  wire        a22_f7_oe,      //       .f7_oe
		input  wire        a22_f0_out,     //       .f0_out
		input  wire        a22_f1_out,     //       .f1_out
		input  wire        a22_f2_out,     //       .f2_out
		input  wire        a22_f3_out,     //       .f3_out
		input  wire        a22_f4_out,     //       .f4_out
		input  wire        a22_f5_out,     //       .f5_out
		input  wire        a22_f6_out,     //       .f6_out
		input  wire        a22_f7_out,     //       .f7_out
		output wire        a22_f_in,       //       .f_in
		inout  wire        a22_GPIO,       //       .GPIO
		input  wire        a23_f0_oe,      //    a23.f0_oe
		input  wire        a23_f1_oe,      //       .f1_oe
		input  wire        a23_f2_oe,      //       .f2_oe
		input  wire        a23_f3_oe,      //       .f3_oe
		input  wire        a23_f4_oe,      //       .f4_oe
		input  wire        a23_f5_oe,      //       .f5_oe
		input  wire        a23_f6_oe,      //       .f6_oe
		input  wire        a23_f7_oe,      //       .f7_oe
		input  wire        a23_f0_out,     //       .f0_out
		input  wire        a23_f1_out,     //       .f1_out
		input  wire        a23_f2_out,     //       .f2_out
		input  wire        a23_f3_out,     //       .f3_out
		input  wire        a23_f4_out,     //       .f4_out
		input  wire        a23_f5_out,     //       .f5_out
		input  wire        a23_f6_out,     //       .f6_out
		input  wire        a23_f7_out,     //       .f7_out
		output wire        a23_f_in,       //       .f_in
		inout  wire        a23_GPIO,       //       .GPIO
		input  wire        a24_f0_oe,      //    a24.f0_oe
		input  wire        a24_f1_oe,      //       .f1_oe
		input  wire        a24_f2_oe,      //       .f2_oe
		input  wire        a24_f3_oe,      //       .f3_oe
		input  wire        a24_f4_oe,      //       .f4_oe
		input  wire        a24_f5_oe,      //       .f5_oe
		input  wire        a24_f6_oe,      //       .f6_oe
		input  wire        a24_f7_oe,      //       .f7_oe
		input  wire        a24_f0_out,     //       .f0_out
		input  wire        a24_f1_out,     //       .f1_out
		input  wire        a24_f2_out,     //       .f2_out
		input  wire        a24_f3_out,     //       .f3_out
		input  wire        a24_f4_out,     //       .f4_out
		input  wire        a24_f5_out,     //       .f5_out
		input  wire        a24_f6_out,     //       .f6_out
		input  wire        a24_f7_out,     //       .f7_out
		output wire        a24_f_in,       //       .f_in
		inout  wire        a24_GPIO,       //       .GPIO
		input  wire        b20_f0_oe,      //    b20.f0_oe
		input  wire        b20_f1_oe,      //       .f1_oe
		input  wire        b20_f2_oe,      //       .f2_oe
		input  wire        b20_f3_oe,      //       .f3_oe
		input  wire        b20_f4_oe,      //       .f4_oe
		input  wire        b20_f5_oe,      //       .f5_oe
		input  wire        b20_f6_oe,      //       .f6_oe
		input  wire        b20_f7_oe,      //       .f7_oe
		input  wire        b20_f0_out,     //       .f0_out
		input  wire        b20_f1_out,     //       .f1_out
		input  wire        b20_f2_out,     //       .f2_out
		input  wire        b20_f3_out,     //       .f3_out
		input  wire        b20_f4_out,     //       .f4_out
		input  wire        b20_f5_out,     //       .f5_out
		input  wire        b20_f6_out,     //       .f6_out
		input  wire        b20_f7_out,     //       .f7_out
		output wire        b20_f_in,       //       .f_in
		inout  wire        b20_GPIO,       //       .GPIO
		input  wire        b21_f0_oe,      //    b21.f0_oe
		input  wire        b21_f1_oe,      //       .f1_oe
		input  wire        b21_f2_oe,      //       .f2_oe
		input  wire        b21_f3_oe,      //       .f3_oe
		input  wire        b21_f4_oe,      //       .f4_oe
		input  wire        b21_f5_oe,      //       .f5_oe
		input  wire        b21_f6_oe,      //       .f6_oe
		input  wire        b21_f7_oe,      //       .f7_oe
		input  wire        b21_f0_out,     //       .f0_out
		input  wire        b21_f1_out,     //       .f1_out
		input  wire        b21_f2_out,     //       .f2_out
		input  wire        b21_f3_out,     //       .f3_out
		input  wire        b21_f4_out,     //       .f4_out
		input  wire        b21_f5_out,     //       .f5_out
		input  wire        b21_f6_out,     //       .f6_out
		input  wire        b21_f7_out,     //       .f7_out
		output wire        b21_f_in,       //       .f_in
		inout  wire        b21_GPIO,       //       .GPIO
		input  wire        b22_f0_oe,      //    b22.f0_oe
		input  wire        b22_f1_oe,      //       .f1_oe
		input  wire        b22_f2_oe,      //       .f2_oe
		input  wire        b22_f3_oe,      //       .f3_oe
		input  wire        b22_f4_oe,      //       .f4_oe
		input  wire        b22_f5_oe,      //       .f5_oe
		input  wire        b22_f6_oe,      //       .f6_oe
		input  wire        b22_f7_oe,      //       .f7_oe
		input  wire        b22_f0_out,     //       .f0_out
		input  wire        b22_f1_out,     //       .f1_out
		input  wire        b22_f2_out,     //       .f2_out
		input  wire        b22_f3_out,     //       .f3_out
		input  wire        b22_f4_out,     //       .f4_out
		input  wire        b22_f5_out,     //       .f5_out
		input  wire        b22_f6_out,     //       .f6_out
		input  wire        b22_f7_out,     //       .f7_out
		output wire        b22_f_in,       //       .f_in
		inout  wire        b22_GPIO,       //       .GPIO
		input  wire        b23_f0_oe,      //    b23.f0_oe
		input  wire        b23_f1_oe,      //       .f1_oe
		input  wire        b23_f2_oe,      //       .f2_oe
		input  wire        b23_f3_oe,      //       .f3_oe
		input  wire        b23_f4_oe,      //       .f4_oe
		input  wire        b23_f5_oe,      //       .f5_oe
		input  wire        b23_f6_oe,      //       .f6_oe
		input  wire        b23_f7_oe,      //       .f7_oe
		input  wire        b23_f0_out,     //       .f0_out
		input  wire        b23_f1_out,     //       .f1_out
		input  wire        b23_f2_out,     //       .f2_out
		input  wire        b23_f3_out,     //       .f3_out
		input  wire        b23_f4_out,     //       .f4_out
		input  wire        b23_f5_out,     //       .f5_out
		input  wire        b23_f6_out,     //       .f6_out
		input  wire        b23_f7_out,     //       .f7_out
		output wire        b23_f_in,       //       .f_in
		inout  wire        b23_GPIO,       //       .GPIO
		input  wire        b24_f0_oe,      //    b24.f0_oe
		input  wire        b24_f1_oe,      //       .f1_oe
		input  wire        b24_f2_oe,      //       .f2_oe
		input  wire        b24_f3_oe,      //       .f3_oe
		input  wire        b24_f4_oe,      //       .f4_oe
		input  wire        b24_f5_oe,      //       .f5_oe
		input  wire        b24_f6_oe,      //       .f6_oe
		input  wire        b24_f7_oe,      //       .f7_oe
		input  wire        b24_f0_out,     //       .f0_out
		input  wire        b24_f1_out,     //       .f1_out
		input  wire        b24_f2_out,     //       .f2_out
		input  wire        b24_f3_out,     //       .f3_out
		input  wire        b24_f4_out,     //       .f4_out
		input  wire        b24_f5_out,     //       .f5_out
		input  wire        b24_f6_out,     //       .f6_out
		input  wire        b24_f7_out,     //       .f7_out
		output wire        b24_f_in,       //       .f_in
		inout  wire        b24_GPIO,       //       .GPIO
		input  wire        shield_A_OCN,   // shield.A_OCN
		output wire        shield_A_PWREN, //       .A_PWREN
		output wire        shield_A_HOE,   //       .A_HOE
		output wire        shield_A_LOE,   //       .A_LOE
		input  wire        shield_B_OCN,   //       .B_OCN
		output wire        shield_B_PWREN, //       .B_PWREN
		output wire        shield_B_HOE,   //       .B_HOE
		output wire        shield_B_LOE,   //       .B_LOE
		input  wire        b25_f0_oe,      //    b25.f0_oe
		input  wire        b25_f1_oe,      //       .f1_oe
		input  wire        b25_f2_oe,      //       .f2_oe
		input  wire        b25_f3_oe,      //       .f3_oe
		input  wire        b25_f4_oe,      //       .f4_oe
		input  wire        b25_f5_oe,      //       .f5_oe
		input  wire        b25_f6_oe,      //       .f6_oe
		input  wire        b25_f7_oe,      //       .f7_oe
		input  wire        b25_f0_out,     //       .f0_out
		input  wire        b25_f1_out,     //       .f1_out
		input  wire        b25_f2_out,     //       .f2_out
		input  wire        b25_f3_out,     //       .f3_out
		input  wire        b25_f4_out,     //       .f4_out
		input  wire        b25_f5_out,     //       .f5_out
		input  wire        b25_f6_out,     //       .f6_out
		input  wire        b25_f7_out,     //       .f7_out
		output wire        b25_f_in,       //       .f_in
		inout  wire        b25_GPIO,       //       .GPIO
		input  wire        a0_f0_oe,       //     a0.f0_oe
		input  wire        a0_f1_oe,       //       .f1_oe
		input  wire        a0_f2_oe,       //       .f2_oe
		input  wire        a0_f3_oe,       //       .f3_oe
		input  wire        a0_f4_oe,       //       .f4_oe
		input  wire        a0_f5_oe,       //       .f5_oe
		input  wire        a0_f6_oe,       //       .f6_oe
		input  wire        a0_f7_oe,       //       .f7_oe
		input  wire        a0_f0_out,      //       .f0_out
		input  wire        a0_f1_out,      //       .f1_out
		input  wire        a0_f2_out,      //       .f2_out
		input  wire        a0_f3_out,      //       .f3_out
		input  wire        a0_f4_out,      //       .f4_out
		input  wire        a0_f5_out,      //       .f5_out
		input  wire        a0_f6_out,      //       .f6_out
		input  wire        a0_f7_out,      //       .f7_out
		output wire        a0_f_in,        //       .f_in
		inout  wire        a0_GPIO,        //       .GPIO
		input  wire        b3_f0_oe,       //     b3.f0_oe
		input  wire        b3_f1_oe,       //       .f1_oe
		input  wire        b3_f2_oe,       //       .f2_oe
		input  wire        b3_f3_oe,       //       .f3_oe
		input  wire        b3_f4_oe,       //       .f4_oe
		input  wire        b3_f5_oe,       //       .f5_oe
		input  wire        b3_f6_oe,       //       .f6_oe
		input  wire        b3_f7_oe,       //       .f7_oe
		input  wire        b3_f0_out,      //       .f0_out
		input  wire        b3_f1_out,      //       .f1_out
		input  wire        b3_f2_out,      //       .f2_out
		input  wire        b3_f3_out,      //       .f3_out
		input  wire        b3_f4_out,      //       .f4_out
		input  wire        b3_f5_out,      //       .f5_out
		input  wire        b3_f6_out,      //       .f6_out
		input  wire        b3_f7_out,      //       .f7_out
		output wire        b3_f_in,        //       .f_in
		inout  wire        b3_GPIO,        //       .GPIO
		input  wire        b2_f0_oe,       //     b2.f0_oe
		input  wire        b2_f1_oe,       //       .f1_oe
		input  wire        b2_f2_oe,       //       .f2_oe
		input  wire        b2_f3_oe,       //       .f3_oe
		input  wire        b2_f4_oe,       //       .f4_oe
		input  wire        b2_f5_oe,       //       .f5_oe
		input  wire        b2_f6_oe,       //       .f6_oe
		input  wire        b2_f7_oe,       //       .f7_oe
		input  wire        b2_f0_out,      //       .f0_out
		input  wire        b2_f1_out,      //       .f1_out
		input  wire        b2_f2_out,      //       .f2_out
		input  wire        b2_f3_out,      //       .f3_out
		input  wire        b2_f4_out,      //       .f4_out
		input  wire        b2_f5_out,      //       .f5_out
		input  wire        b2_f6_out,      //       .f6_out
		input  wire        b2_f7_out,      //       .f7_out
		output wire        b2_f_in,        //       .f_in
		inout  wire        b2_GPIO,        //       .GPIO
		output wire        led_f0_R,       // led_f0.R
		output wire        led_f0_G,       //       .G
		output wire        led_f0_B,       //       .B
		input  wire        b5_f0_oe,       //     b5.f0_oe
		input  wire        b5_f1_oe,       //       .f1_oe
		input  wire        b5_f2_oe,       //       .f2_oe
		input  wire        b5_f3_oe,       //       .f3_oe
		input  wire        b5_f4_oe,       //       .f4_oe
		input  wire        b5_f5_oe,       //       .f5_oe
		input  wire        b5_f6_oe,       //       .f6_oe
		input  wire        b5_f7_oe,       //       .f7_oe
		input  wire        b5_f0_out,      //       .f0_out
		input  wire        b5_f1_out,      //       .f1_out
		input  wire        b5_f2_out,      //       .f2_out
		input  wire        b5_f3_out,      //       .f3_out
		input  wire        b5_f4_out,      //       .f4_out
		input  wire        b5_f5_out,      //       .f5_out
		input  wire        b5_f6_out,      //       .f6_out
		input  wire        b5_f7_out,      //       .f7_out
		output wire        b5_f_in,        //       .f_in
		inout  wire        b5_GPIO,        //       .GPIO
		output wire        led_f1_R,       // led_f1.R
		output wire        led_f1_G,       //       .G
		output wire        led_f1_B,       //       .B
		input  wire        b4_f0_oe,       //     b4.f0_oe
		input  wire        b4_f1_oe,       //       .f1_oe
		input  wire        b4_f2_oe,       //       .f2_oe
		input  wire        b4_f3_oe,       //       .f3_oe
		input  wire        b4_f4_oe,       //       .f4_oe
		input  wire        b4_f5_oe,       //       .f5_oe
		input  wire        b4_f6_oe,       //       .f6_oe
		input  wire        b4_f7_oe,       //       .f7_oe
		input  wire        b4_f0_out,      //       .f0_out
		input  wire        b4_f1_out,      //       .f1_out
		input  wire        b4_f2_out,      //       .f2_out
		input  wire        b4_f3_out,      //       .f3_out
		input  wire        b4_f4_out,      //       .f4_out
		input  wire        b4_f5_out,      //       .f5_out
		input  wire        b4_f6_out,      //       .f6_out
		input  wire        b4_f7_out,      //       .f7_out
		output wire        b4_f_in,        //       .f_in
		inout  wire        b4_GPIO,        //       .GPIO
		input  wire        b7_f0_oe,       //     b7.f0_oe
		input  wire        b7_f1_oe,       //       .f1_oe
		input  wire        b7_f2_oe,       //       .f2_oe
		input  wire        b7_f3_oe,       //       .f3_oe
		input  wire        b7_f4_oe,       //       .f4_oe
		input  wire        b7_f5_oe,       //       .f5_oe
		input  wire        b7_f6_oe,       //       .f6_oe
		input  wire        b7_f7_oe,       //       .f7_oe
		input  wire        b7_f0_out,      //       .f0_out
		input  wire        b7_f1_out,      //       .f1_out
		input  wire        b7_f2_out,      //       .f2_out
		input  wire        b7_f3_out,      //       .f3_out
		input  wire        b7_f4_out,      //       .f4_out
		input  wire        b7_f5_out,      //       .f5_out
		input  wire        b7_f6_out,      //       .f6_out
		input  wire        b7_f7_out,      //       .f7_out
		output wire        b7_f_in,        //       .f_in
		inout  wire        b7_GPIO,        //       .GPIO
		input  wire        b6_f0_oe,       //     b6.f0_oe
		input  wire        b6_f1_oe,       //       .f1_oe
		input  wire        b6_f2_oe,       //       .f2_oe
		input  wire        b6_f3_oe,       //       .f3_oe
		input  wire        b6_f4_oe,       //       .f4_oe
		input  wire        b6_f5_oe,       //       .f5_oe
		input  wire        b6_f6_oe,       //       .f6_oe
		input  wire        b6_f7_oe,       //       .f7_oe
		input  wire        b6_f0_out,      //       .f0_out
		input  wire        b6_f1_out,      //       .f1_out
		input  wire        b6_f2_out,      //       .f2_out
		input  wire        b6_f3_out,      //       .f3_out
		input  wire        b6_f4_out,      //       .f4_out
		input  wire        b6_f5_out,      //       .f5_out
		input  wire        b6_f6_out,      //       .f6_out
		input  wire        b6_f7_out,      //       .f7_out
		output wire        b6_f_in,        //       .f_in
		inout  wire        b6_GPIO,        //       .GPIO
		input  wire        b9_f0_oe,       //     b9.f0_oe
		input  wire        b9_f1_oe,       //       .f1_oe
		input  wire        b9_f2_oe,       //       .f2_oe
		input  wire        b9_f3_oe,       //       .f3_oe
		input  wire        b9_f4_oe,       //       .f4_oe
		input  wire        b9_f5_oe,       //       .f5_oe
		input  wire        b9_f6_oe,       //       .f6_oe
		input  wire        b9_f7_oe,       //       .f7_oe
		input  wire        b9_f0_out,      //       .f0_out
		input  wire        b9_f1_out,      //       .f1_out
		input  wire        b9_f2_out,      //       .f2_out
		input  wire        b9_f3_out,      //       .f3_out
		input  wire        b9_f4_out,      //       .f4_out
		input  wire        b9_f5_out,      //       .f5_out
		input  wire        b9_f6_out,      //       .f6_out
		input  wire        b9_f7_out,      //       .f7_out
		output wire        b9_f_in,        //       .f_in
		inout  wire        b9_GPIO,        //       .GPIO
		input  wire        b8_f0_oe,       //     b8.f0_oe
		input  wire        b8_f1_oe,       //       .f1_oe
		input  wire        b8_f2_oe,       //       .f2_oe
		input  wire        b8_f3_oe,       //       .f3_oe
		input  wire        b8_f4_oe,       //       .f4_oe
		input  wire        b8_f5_oe,       //       .f5_oe
		input  wire        b8_f6_oe,       //       .f6_oe
		input  wire        b8_f7_oe,       //       .f7_oe
		input  wire        b8_f0_out,      //       .f0_out
		input  wire        b8_f1_out,      //       .f1_out
		input  wire        b8_f2_out,      //       .f2_out
		input  wire        b8_f3_out,      //       .f3_out
		input  wire        b8_f4_out,      //       .f4_out
		input  wire        b8_f5_out,      //       .f5_out
		input  wire        b8_f6_out,      //       .f6_out
		input  wire        b8_f7_out,      //       .f7_out
		output wire        b8_f_in,        //       .f_in
		inout  wire        b8_GPIO,        //       .GPIO
		input  wire        a9_f0_oe,       //     a9.f0_oe
		input  wire        a9_f1_oe,       //       .f1_oe
		input  wire        a9_f2_oe,       //       .f2_oe
		input  wire        a9_f3_oe,       //       .f3_oe
		input  wire        a9_f4_oe,       //       .f4_oe
		input  wire        a9_f5_oe,       //       .f5_oe
		input  wire        a9_f6_oe,       //       .f6_oe
		input  wire        a9_f7_oe,       //       .f7_oe
		input  wire        a9_f0_out,      //       .f0_out
		input  wire        a9_f1_out,      //       .f1_out
		input  wire        a9_f2_out,      //       .f2_out
		input  wire        a9_f3_out,      //       .f3_out
		input  wire        a9_f4_out,      //       .f4_out
		input  wire        a9_f5_out,      //       .f5_out
		input  wire        a9_f6_out,      //       .f6_out
		input  wire        a9_f7_out,      //       .f7_out
		output wire        a9_f_in,        //       .f_in
		inout  wire        a9_GPIO,        //       .GPIO
		input  wire        b0_f0_oe,       //     b0.f0_oe
		input  wire        b0_f1_oe,       //       .f1_oe
		input  wire        b0_f2_oe,       //       .f2_oe
		input  wire        b0_f3_oe,       //       .f3_oe
		input  wire        b0_f4_oe,       //       .f4_oe
		input  wire        b0_f5_oe,       //       .f5_oe
		input  wire        b0_f6_oe,       //       .f6_oe
		input  wire        b0_f7_oe,       //       .f7_oe
		input  wire        b0_f0_out,      //       .f0_out
		input  wire        b0_f1_out,      //       .f1_out
		input  wire        b0_f2_out,      //       .f2_out
		input  wire        b0_f3_out,      //       .f3_out
		input  wire        b0_f4_out,      //       .f4_out
		input  wire        b0_f5_out,      //       .f5_out
		input  wire        b0_f6_out,      //       .f6_out
		input  wire        b0_f7_out,      //       .f7_out
		output wire        b0_f_in,        //       .f_in
		inout  wire        b0_GPIO,        //       .GPIO
		input  wire        b1_f0_oe,       //     b1.f0_oe
		input  wire        b1_f1_oe,       //       .f1_oe
		input  wire        b1_f2_oe,       //       .f2_oe
		input  wire        b1_f3_oe,       //       .f3_oe
		input  wire        b1_f4_oe,       //       .f4_oe
		input  wire        b1_f5_oe,       //       .f5_oe
		input  wire        b1_f6_oe,       //       .f6_oe
		input  wire        b1_f7_oe,       //       .f7_oe
		input  wire        b1_f0_out,      //       .f0_out
		input  wire        b1_f1_out,      //       .f1_out
		input  wire        b1_f2_out,      //       .f2_out
		input  wire        b1_f3_out,      //       .f3_out
		input  wire        b1_f4_out,      //       .f4_out
		input  wire        b1_f5_out,      //       .f5_out
		input  wire        b1_f6_out,      //       .f6_out
		input  wire        b1_f7_out,      //       .f7_out
		output wire        b1_f_in,        //       .f_in
		inout  wire        b1_GPIO,        //       .GPIO
		input  wire        a1_f0_oe,       //     a1.f0_oe
		input  wire        a1_f1_oe,       //       .f1_oe
		input  wire        a1_f2_oe,       //       .f2_oe
		input  wire        a1_f3_oe,       //       .f3_oe
		input  wire        a1_f4_oe,       //       .f4_oe
		input  wire        a1_f5_oe,       //       .f5_oe
		input  wire        a1_f6_oe,       //       .f6_oe
		input  wire        a1_f7_oe,       //       .f7_oe
		input  wire        a1_f0_out,      //       .f0_out
		input  wire        a1_f1_out,      //       .f1_out
		input  wire        a1_f2_out,      //       .f2_out
		input  wire        a1_f3_out,      //       .f3_out
		input  wire        a1_f4_out,      //       .f4_out
		input  wire        a1_f5_out,      //       .f5_out
		input  wire        a1_f6_out,      //       .f6_out
		input  wire        a1_f7_out,      //       .f7_out
		output wire        a1_f_in,        //       .f_in
		inout  wire        a1_GPIO,        //       .GPIO
		input  wire        a2_f0_oe,       //     a2.f0_oe
		input  wire        a2_f1_oe,       //       .f1_oe
		input  wire        a2_f2_oe,       //       .f2_oe
		input  wire        a2_f3_oe,       //       .f3_oe
		input  wire        a2_f4_oe,       //       .f4_oe
		input  wire        a2_f5_oe,       //       .f5_oe
		input  wire        a2_f6_oe,       //       .f6_oe
		input  wire        a2_f7_oe,       //       .f7_oe
		input  wire        a2_f0_out,      //       .f0_out
		input  wire        a2_f1_out,      //       .f1_out
		input  wire        a2_f2_out,      //       .f2_out
		input  wire        a2_f3_out,      //       .f3_out
		input  wire        a2_f4_out,      //       .f4_out
		input  wire        a2_f5_out,      //       .f5_out
		input  wire        a2_f6_out,      //       .f6_out
		input  wire        a2_f7_out,      //       .f7_out
		output wire        a2_f_in,        //       .f_in
		inout  wire        a2_GPIO,        //       .GPIO
		input  wire        a3_f0_oe,       //     a3.f0_oe
		input  wire        a3_f1_oe,       //       .f1_oe
		input  wire        a3_f2_oe,       //       .f2_oe
		input  wire        a3_f3_oe,       //       .f3_oe
		input  wire        a3_f4_oe,       //       .f4_oe
		input  wire        a3_f5_oe,       //       .f5_oe
		input  wire        a3_f6_oe,       //       .f6_oe
		input  wire        a3_f7_oe,       //       .f7_oe
		input  wire        a3_f0_out,      //       .f0_out
		input  wire        a3_f1_out,      //       .f1_out
		input  wire        a3_f2_out,      //       .f2_out
		input  wire        a3_f3_out,      //       .f3_out
		input  wire        a3_f4_out,      //       .f4_out
		input  wire        a3_f5_out,      //       .f5_out
		input  wire        a3_f6_out,      //       .f6_out
		input  wire        a3_f7_out,      //       .f7_out
		output wire        a3_f_in,        //       .f_in
		inout  wire        a3_GPIO,        //       .GPIO
		input  wire        a4_f0_oe,       //     a4.f0_oe
		input  wire        a4_f1_oe,       //       .f1_oe
		input  wire        a4_f2_oe,       //       .f2_oe
		input  wire        a4_f3_oe,       //       .f3_oe
		input  wire        a4_f4_oe,       //       .f4_oe
		input  wire        a4_f5_oe,       //       .f5_oe
		input  wire        a4_f6_oe,       //       .f6_oe
		input  wire        a4_f7_oe,       //       .f7_oe
		input  wire        a4_f0_out,      //       .f0_out
		input  wire        a4_f1_out,      //       .f1_out
		input  wire        a4_f2_out,      //       .f2_out
		input  wire        a4_f3_out,      //       .f3_out
		input  wire        a4_f4_out,      //       .f4_out
		input  wire        a4_f5_out,      //       .f5_out
		input  wire        a4_f6_out,      //       .f6_out
		input  wire        a4_f7_out,      //       .f7_out
		output wire        a4_f_in,        //       .f_in
		inout  wire        a4_GPIO,        //       .GPIO
		input  wire        a5_f0_oe,       //     a5.f0_oe
		input  wire        a5_f1_oe,       //       .f1_oe
		input  wire        a5_f2_oe,       //       .f2_oe
		input  wire        a5_f3_oe,       //       .f3_oe
		input  wire        a5_f4_oe,       //       .f4_oe
		input  wire        a5_f5_oe,       //       .f5_oe
		input  wire        a5_f6_oe,       //       .f6_oe
		input  wire        a5_f7_oe,       //       .f7_oe
		input  wire        a5_f0_out,      //       .f0_out
		input  wire        a5_f1_out,      //       .f1_out
		input  wire        a5_f2_out,      //       .f2_out
		input  wire        a5_f3_out,      //       .f3_out
		input  wire        a5_f4_out,      //       .f4_out
		input  wire        a5_f5_out,      //       .f5_out
		input  wire        a5_f6_out,      //       .f6_out
		input  wire        a5_f7_out,      //       .f7_out
		output wire        a5_f_in,        //       .f_in
		inout  wire        a5_GPIO,        //       .GPIO
		input  wire        a6_f0_oe,       //     a6.f0_oe
		input  wire        a6_f1_oe,       //       .f1_oe
		input  wire        a6_f2_oe,       //       .f2_oe
		input  wire        a6_f3_oe,       //       .f3_oe
		input  wire        a6_f4_oe,       //       .f4_oe
		input  wire        a6_f5_oe,       //       .f5_oe
		input  wire        a6_f6_oe,       //       .f6_oe
		input  wire        a6_f7_oe,       //       .f7_oe
		input  wire        a6_f0_out,      //       .f0_out
		input  wire        a6_f1_out,      //       .f1_out
		input  wire        a6_f2_out,      //       .f2_out
		input  wire        a6_f3_out,      //       .f3_out
		input  wire        a6_f4_out,      //       .f4_out
		input  wire        a6_f5_out,      //       .f5_out
		input  wire        a6_f6_out,      //       .f6_out
		input  wire        a6_f7_out,      //       .f7_out
		output wire        a6_f_in,        //       .f_in
		inout  wire        a6_GPIO,        //       .GPIO
		input  wire        a7_f0_oe,       //     a7.f0_oe
		input  wire        a7_f1_oe,       //       .f1_oe
		input  wire        a7_f2_oe,       //       .f2_oe
		input  wire        a7_f3_oe,       //       .f3_oe
		input  wire        a7_f4_oe,       //       .f4_oe
		input  wire        a7_f5_oe,       //       .f5_oe
		input  wire        a7_f6_oe,       //       .f6_oe
		input  wire        a7_f7_oe,       //       .f7_oe
		input  wire        a7_f0_out,      //       .f0_out
		input  wire        a7_f1_out,      //       .f1_out
		input  wire        a7_f2_out,      //       .f2_out
		input  wire        a7_f3_out,      //       .f3_out
		input  wire        a7_f4_out,      //       .f4_out
		input  wire        a7_f5_out,      //       .f5_out
		input  wire        a7_f6_out,      //       .f6_out
		input  wire        a7_f7_out,      //       .f7_out
		output wire        a7_f_in,        //       .f_in
		inout  wire        a7_GPIO,        //       .GPIO
		input  wire        a8_f0_oe,       //     a8.f0_oe
		input  wire        a8_f1_oe,       //       .f1_oe
		input  wire        a8_f2_oe,       //       .f2_oe
		input  wire        a8_f3_oe,       //       .f3_oe
		input  wire        a8_f4_oe,       //       .f4_oe
		input  wire        a8_f5_oe,       //       .f5_oe
		input  wire        a8_f6_oe,       //       .f6_oe
		input  wire        a8_f7_oe,       //       .f7_oe
		input  wire        a8_f0_out,      //       .f0_out
		input  wire        a8_f1_out,      //       .f1_out
		input  wire        a8_f2_out,      //       .f2_out
		input  wire        a8_f3_out,      //       .f3_out
		input  wire        a8_f4_out,      //       .f4_out
		input  wire        a8_f5_out,      //       .f5_out
		input  wire        a8_f6_out,      //       .f6_out
		input  wire        a8_f7_out,      //       .f7_out
		output wire        a8_f_in,        //       .f_in
		inout  wire        a8_GPIO         //       .GPIO
	);

	wire         sam9_mrst_reset;                                                                         // SAM9:rso_MRST_reset -> [FuncLED_0:rsi_MRST_reset, FuncLED_0_LEDD_translator:reset, FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:reset, FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FuncLED_1:rsi_MRST_reset, FuncLED_1_LEDD_translator:reset, FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:reset, FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FuncLED_2:rsi_MRST_reset, FuncLED_2_LEDD_translator:reset, FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:reset, FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FuncLED_3:rsi_MRST_reset, FuncLED_3_LEDD_translator:reset, FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:reset, FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SAM9_M1_translator:reset, SAM9_M1_translator_avalon_universal_master_0_agent:reset, Shield_Admin:rsi_MRST_reset, Shield_Admin_Ctrl_translator:reset, Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:reset, Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A0:rsi_MRST_reset, Shiled_IO_A0_ctrl_translator:reset, Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A10:rsi_MRST_reset, Shiled_IO_A10_ctrl_translator:reset, Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A11:rsi_MRST_reset, Shiled_IO_A11_ctrl_translator:reset, Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A12:rsi_MRST_reset, Shiled_IO_A12_ctrl_translator:reset, Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A13:rsi_MRST_reset, Shiled_IO_A13_ctrl_translator:reset, Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A14:rsi_MRST_reset, Shiled_IO_A14_ctrl_translator:reset, Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A15:rsi_MRST_reset, Shiled_IO_A15_ctrl_translator:reset, Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A16:rsi_MRST_reset, Shiled_IO_A16_ctrl_translator:reset, Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A17:rsi_MRST_reset, Shiled_IO_A17_ctrl_translator:reset, Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A18:rsi_MRST_reset, Shiled_IO_A18_ctrl_translator:reset, Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A19:rsi_MRST_reset, Shiled_IO_A19_ctrl_translator:reset, Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A1:rsi_MRST_reset, Shiled_IO_A1_ctrl_translator:reset, Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A20:rsi_MRST_reset, Shiled_IO_A20_ctrl_translator:reset, Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A21:rsi_MRST_reset, Shiled_IO_A21_ctrl_translator:reset, Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A22:rsi_MRST_reset, Shiled_IO_A22_ctrl_translator:reset, Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A23:rsi_MRST_reset, Shiled_IO_A23_ctrl_translator:reset, Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A24:rsi_MRST_reset, Shiled_IO_A24_ctrl_translator:reset, Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A25:rsi_MRST_reset, Shiled_IO_A25_ctrl_translator:reset, Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A2:rsi_MRST_reset, Shiled_IO_A2_ctrl_translator:reset, Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A3:rsi_MRST_reset, Shiled_IO_A3_ctrl_translator:reset, Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A4:rsi_MRST_reset, Shiled_IO_A4_ctrl_translator:reset, Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A5:rsi_MRST_reset, Shiled_IO_A5_ctrl_translator:reset, Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A6:rsi_MRST_reset, Shiled_IO_A6_ctrl_translator:reset, Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A7:rsi_MRST_reset, Shiled_IO_A7_ctrl_translator:reset, Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A8:rsi_MRST_reset, Shiled_IO_A8_ctrl_translator:reset, Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_A9:rsi_MRST_reset, Shiled_IO_A9_ctrl_translator:reset, Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B0:rsi_MRST_reset, Shiled_IO_B0_ctrl_translator:reset, Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B10:rsi_MRST_reset, Shiled_IO_B10_ctrl_translator:reset, Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B11:rsi_MRST_reset, Shiled_IO_B11_ctrl_translator:reset, Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B12:rsi_MRST_reset, Shiled_IO_B12_ctrl_translator:reset, Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B13:rsi_MRST_reset, Shiled_IO_B13_ctrl_translator:reset, Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B14:rsi_MRST_reset, Shiled_IO_B14_ctrl_translator:reset, Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B15:rsi_MRST_reset, Shiled_IO_B15_ctrl_translator:reset, Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B16:rsi_MRST_reset, Shiled_IO_B16_ctrl_translator:reset, Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B17:rsi_MRST_reset, Shiled_IO_B17_ctrl_translator:reset, Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B18:rsi_MRST_reset, Shiled_IO_B18_ctrl_translator:reset, Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B19:rsi_MRST_reset, Shiled_IO_B19_ctrl_translator:reset, Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B1:rsi_MRST_reset, Shiled_IO_B1_ctrl_translator:reset, Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B20:rsi_MRST_reset, Shiled_IO_B20_ctrl_translator:reset, Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B21:rsi_MRST_reset, Shiled_IO_B21_ctrl_translator:reset, Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B22:rsi_MRST_reset, Shiled_IO_B22_ctrl_translator:reset, Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B23:rsi_MRST_reset, Shiled_IO_B23_ctrl_translator:reset, Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B24:rsi_MRST_reset, Shiled_IO_B24_ctrl_translator:reset, Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B25:rsi_MRST_reset, Shiled_IO_B25_ctrl_translator:reset, Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B2:rsi_MRST_reset, Shiled_IO_B2_ctrl_translator:reset, Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B3:rsi_MRST_reset, Shiled_IO_B3_ctrl_translator:reset, Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B4:rsi_MRST_reset, Shiled_IO_B4_ctrl_translator:reset, Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B5:rsi_MRST_reset, Shiled_IO_B5_ctrl_translator:reset, Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B6:rsi_MRST_reset, Shiled_IO_B6_ctrl_translator:reset, Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B7:rsi_MRST_reset, Shiled_IO_B7_ctrl_translator:reset, Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B8:rsi_MRST_reset, Shiled_IO_B8_ctrl_translator:reset, Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shiled_IO_B9:rsi_MRST_reset, Shiled_IO_B9_ctrl_translator:reset, Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:reset, Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SysID:rsi_MRST_reset, SysID_SysID_translator:reset, SysID_SysID_translator_avalon_universal_slave_0_agent:reset, SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, burst_adapter_004:reset, burst_adapter_005:reset, burst_adapter_006:reset, burst_adapter_007:reset, burst_adapter_008:reset, burst_adapter_009:reset, burst_adapter_010:reset, burst_adapter_011:reset, burst_adapter_012:reset, burst_adapter_013:reset, burst_adapter_014:reset, burst_adapter_015:reset, burst_adapter_016:reset, burst_adapter_017:reset, burst_adapter_018:reset, burst_adapter_019:reset, burst_adapter_020:reset, burst_adapter_021:reset, burst_adapter_022:reset, burst_adapter_023:reset, burst_adapter_024:reset, burst_adapter_025:reset, burst_adapter_026:reset, burst_adapter_027:reset, burst_adapter_028:reset, burst_adapter_029:reset, burst_adapter_030:reset, burst_adapter_031:reset, burst_adapter_032:reset, burst_adapter_033:reset, burst_adapter_034:reset, burst_adapter_035:reset, burst_adapter_036:reset, burst_adapter_037:reset, burst_adapter_038:reset, burst_adapter_039:reset, burst_adapter_040:reset, burst_adapter_041:reset, burst_adapter_042:reset, burst_adapter_043:reset, burst_adapter_044:reset, burst_adapter_045:reset, burst_adapter_046:reset, burst_adapter_047:reset, burst_adapter_048:reset, burst_adapter_049:reset, burst_adapter_050:reset, burst_adapter_051:reset, cmd_xbar_demux:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, id_router_025:reset, id_router_026:reset, id_router_027:reset, id_router_028:reset, id_router_029:reset, id_router_030:reset, id_router_031:reset, id_router_032:reset, id_router_033:reset, id_router_034:reset, id_router_035:reset, id_router_036:reset, id_router_037:reset, id_router_038:reset, id_router_039:reset, id_router_040:reset, id_router_041:reset, id_router_042:reset, id_router_043:reset, id_router_044:reset, id_router_045:reset, id_router_046:reset, id_router_047:reset, id_router_048:reset, id_router_049:reset, id_router_050:reset, id_router_051:reset, id_router_052:reset, id_router_053:reset, id_router_054:reset, id_router_055:reset, id_router_056:reset, id_router_057:reset, irq_mapper:reset, irq_synchronizer:receiver_reset, irq_synchronizer:sender_reset, limiter:reset, qsys_test_LEDState_0:rsi_MRST_reset, qsys_test_LEDState_1:rsi_MRST_reset, qsys_test_LEDState_2:rsi_MRST_reset, qsys_test_LEDState_3:rsi_MRST_reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, rsp_xbar_demux_025:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, rsp_xbar_demux_029:reset, rsp_xbar_demux_030:reset, rsp_xbar_demux_031:reset, rsp_xbar_demux_032:reset, rsp_xbar_demux_033:reset, rsp_xbar_demux_034:reset, rsp_xbar_demux_035:reset, rsp_xbar_demux_036:reset, rsp_xbar_demux_037:reset, rsp_xbar_demux_038:reset, rsp_xbar_demux_039:reset, rsp_xbar_demux_040:reset, rsp_xbar_demux_041:reset, rsp_xbar_demux_042:reset, rsp_xbar_demux_043:reset, rsp_xbar_demux_044:reset, rsp_xbar_demux_045:reset, rsp_xbar_demux_046:reset, rsp_xbar_demux_047:reset, rsp_xbar_demux_048:reset, rsp_xbar_demux_049:reset, rsp_xbar_demux_050:reset, rsp_xbar_demux_051:reset, rsp_xbar_demux_052:reset, rsp_xbar_demux_053:reset, rsp_xbar_demux_054:reset, rsp_xbar_demux_055:reset, rsp_xbar_demux_056:reset, rsp_xbar_demux_057:reset, rsp_xbar_mux:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset, width_adapter_008:reset, width_adapter_009:reset, width_adapter_010:reset, width_adapter_011:reset, width_adapter_012:reset, width_adapter_013:reset, width_adapter_014:reset, width_adapter_015:reset, width_adapter_016:reset, width_adapter_017:reset, width_adapter_018:reset, width_adapter_019:reset, width_adapter_020:reset, width_adapter_021:reset, width_adapter_022:reset, width_adapter_023:reset, width_adapter_024:reset, width_adapter_025:reset, width_adapter_026:reset, width_adapter_027:reset, width_adapter_028:reset, width_adapter_029:reset, width_adapter_030:reset, width_adapter_031:reset, width_adapter_032:reset, width_adapter_033:reset, width_adapter_034:reset, width_adapter_035:reset, width_adapter_036:reset, width_adapter_037:reset, width_adapter_038:reset, width_adapter_039:reset, width_adapter_040:reset, width_adapter_041:reset, width_adapter_042:reset, width_adapter_043:reset, width_adapter_044:reset, width_adapter_045:reset, width_adapter_046:reset, width_adapter_047:reset, width_adapter_048:reset, width_adapter_049:reset, width_adapter_050:reset, width_adapter_051:reset, width_adapter_052:reset, width_adapter_053:reset, width_adapter_054:reset, width_adapter_055:reset, width_adapter_056:reset, width_adapter_057:reset, width_adapter_058:reset, width_adapter_059:reset, width_adapter_060:reset, width_adapter_061:reset, width_adapter_062:reset, width_adapter_063:reset, width_adapter_064:reset, width_adapter_065:reset, width_adapter_066:reset, width_adapter_067:reset, width_adapter_068:reset, width_adapter_069:reset, width_adapter_070:reset, width_adapter_071:reset, width_adapter_072:reset, width_adapter_073:reset, width_adapter_074:reset, width_adapter_075:reset, width_adapter_076:reset, width_adapter_077:reset, width_adapter_078:reset, width_adapter_079:reset, width_adapter_080:reset, width_adapter_081:reset, width_adapter_082:reset, width_adapter_083:reset, width_adapter_084:reset, width_adapter_085:reset, width_adapter_086:reset, width_adapter_087:reset, width_adapter_088:reset, width_adapter_089:reset, width_adapter_090:reset, width_adapter_091:reset, width_adapter_092:reset, width_adapter_093:reset, width_adapter_094:reset, width_adapter_095:reset, width_adapter_096:reset, width_adapter_097:reset, width_adapter_098:reset, width_adapter_099:reset, width_adapter_100:reset, width_adapter_101:reset, width_adapter_102:reset, width_adapter_103:reset]
	wire         sam9_mclk_clk;                                                                           // SAM9:cso_MCLK_clk -> [FuncLED_0:csi_MCLK_clk, FuncLED_0_LEDD_translator:clk, FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:clk, FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, FuncLED_1:csi_MCLK_clk, FuncLED_1_LEDD_translator:clk, FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:clk, FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, FuncLED_2:csi_MCLK_clk, FuncLED_2_LEDD_translator:clk, FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:clk, FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, FuncLED_3:csi_MCLK_clk, FuncLED_3_LEDD_translator:clk, FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:clk, FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, SAM9_M1_translator:clk, SAM9_M1_translator_avalon_universal_master_0_agent:clk, Shield_Admin:csi_MCLK_clk, Shield_Admin_Ctrl_translator:clk, Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:clk, Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A0:csi_MCLK_clk, Shiled_IO_A0_ctrl_translator:clk, Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A10:csi_MCLK_clk, Shiled_IO_A10_ctrl_translator:clk, Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A11:csi_MCLK_clk, Shiled_IO_A11_ctrl_translator:clk, Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A12:csi_MCLK_clk, Shiled_IO_A12_ctrl_translator:clk, Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A13:csi_MCLK_clk, Shiled_IO_A13_ctrl_translator:clk, Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A14:csi_MCLK_clk, Shiled_IO_A14_ctrl_translator:clk, Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A15:csi_MCLK_clk, Shiled_IO_A15_ctrl_translator:clk, Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A16:csi_MCLK_clk, Shiled_IO_A16_ctrl_translator:clk, Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A17:csi_MCLK_clk, Shiled_IO_A17_ctrl_translator:clk, Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A18:csi_MCLK_clk, Shiled_IO_A18_ctrl_translator:clk, Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A19:csi_MCLK_clk, Shiled_IO_A19_ctrl_translator:clk, Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A1:csi_MCLK_clk, Shiled_IO_A1_ctrl_translator:clk, Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A20:csi_MCLK_clk, Shiled_IO_A20_ctrl_translator:clk, Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A21:csi_MCLK_clk, Shiled_IO_A21_ctrl_translator:clk, Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A22:csi_MCLK_clk, Shiled_IO_A22_ctrl_translator:clk, Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A23:csi_MCLK_clk, Shiled_IO_A23_ctrl_translator:clk, Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A24:csi_MCLK_clk, Shiled_IO_A24_ctrl_translator:clk, Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A25:csi_MCLK_clk, Shiled_IO_A25_ctrl_translator:clk, Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A2:csi_MCLK_clk, Shiled_IO_A2_ctrl_translator:clk, Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A3:csi_MCLK_clk, Shiled_IO_A3_ctrl_translator:clk, Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A4:csi_MCLK_clk, Shiled_IO_A4_ctrl_translator:clk, Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A5:csi_MCLK_clk, Shiled_IO_A5_ctrl_translator:clk, Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A6:csi_MCLK_clk, Shiled_IO_A6_ctrl_translator:clk, Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A7:csi_MCLK_clk, Shiled_IO_A7_ctrl_translator:clk, Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A8:csi_MCLK_clk, Shiled_IO_A8_ctrl_translator:clk, Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_A9:csi_MCLK_clk, Shiled_IO_A9_ctrl_translator:clk, Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B0:csi_MCLK_clk, Shiled_IO_B0_ctrl_translator:clk, Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B10:csi_MCLK_clk, Shiled_IO_B10_ctrl_translator:clk, Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B11:csi_MCLK_clk, Shiled_IO_B11_ctrl_translator:clk, Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B12:csi_MCLK_clk, Shiled_IO_B12_ctrl_translator:clk, Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B13:csi_MCLK_clk, Shiled_IO_B13_ctrl_translator:clk, Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B14:csi_MCLK_clk, Shiled_IO_B14_ctrl_translator:clk, Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B15:csi_MCLK_clk, Shiled_IO_B15_ctrl_translator:clk, Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B16:csi_MCLK_clk, Shiled_IO_B16_ctrl_translator:clk, Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B17:csi_MCLK_clk, Shiled_IO_B17_ctrl_translator:clk, Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B18:csi_MCLK_clk, Shiled_IO_B18_ctrl_translator:clk, Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B19:csi_MCLK_clk, Shiled_IO_B19_ctrl_translator:clk, Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B1:csi_MCLK_clk, Shiled_IO_B1_ctrl_translator:clk, Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B20:csi_MCLK_clk, Shiled_IO_B20_ctrl_translator:clk, Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B21:csi_MCLK_clk, Shiled_IO_B21_ctrl_translator:clk, Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B22:csi_MCLK_clk, Shiled_IO_B22_ctrl_translator:clk, Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B23:csi_MCLK_clk, Shiled_IO_B23_ctrl_translator:clk, Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B24:csi_MCLK_clk, Shiled_IO_B24_ctrl_translator:clk, Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B25:csi_MCLK_clk, Shiled_IO_B25_ctrl_translator:clk, Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B2:csi_MCLK_clk, Shiled_IO_B2_ctrl_translator:clk, Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B3:csi_MCLK_clk, Shiled_IO_B3_ctrl_translator:clk, Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B4:csi_MCLK_clk, Shiled_IO_B4_ctrl_translator:clk, Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B5:csi_MCLK_clk, Shiled_IO_B5_ctrl_translator:clk, Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B6:csi_MCLK_clk, Shiled_IO_B6_ctrl_translator:clk, Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B7:csi_MCLK_clk, Shiled_IO_B7_ctrl_translator:clk, Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B8:csi_MCLK_clk, Shiled_IO_B8_ctrl_translator:clk, Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shiled_IO_B9:csi_MCLK_clk, Shiled_IO_B9_ctrl_translator:clk, Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:clk, Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, SysID:csi_MCLK_clk, SysID_SysID_translator:clk, SysID_SysID_translator_avalon_universal_slave_0_agent:clk, SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, burst_adapter_003:clk, burst_adapter_004:clk, burst_adapter_005:clk, burst_adapter_006:clk, burst_adapter_007:clk, burst_adapter_008:clk, burst_adapter_009:clk, burst_adapter_010:clk, burst_adapter_011:clk, burst_adapter_012:clk, burst_adapter_013:clk, burst_adapter_014:clk, burst_adapter_015:clk, burst_adapter_016:clk, burst_adapter_017:clk, burst_adapter_018:clk, burst_adapter_019:clk, burst_adapter_020:clk, burst_adapter_021:clk, burst_adapter_022:clk, burst_adapter_023:clk, burst_adapter_024:clk, burst_adapter_025:clk, burst_adapter_026:clk, burst_adapter_027:clk, burst_adapter_028:clk, burst_adapter_029:clk, burst_adapter_030:clk, burst_adapter_031:clk, burst_adapter_032:clk, burst_adapter_033:clk, burst_adapter_034:clk, burst_adapter_035:clk, burst_adapter_036:clk, burst_adapter_037:clk, burst_adapter_038:clk, burst_adapter_039:clk, burst_adapter_040:clk, burst_adapter_041:clk, burst_adapter_042:clk, burst_adapter_043:clk, burst_adapter_044:clk, burst_adapter_045:clk, burst_adapter_046:clk, burst_adapter_047:clk, burst_adapter_048:clk, burst_adapter_049:clk, burst_adapter_050:clk, burst_adapter_051:clk, cmd_xbar_demux:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, id_router_019:clk, id_router_020:clk, id_router_021:clk, id_router_022:clk, id_router_023:clk, id_router_024:clk, id_router_025:clk, id_router_026:clk, id_router_027:clk, id_router_028:clk, id_router_029:clk, id_router_030:clk, id_router_031:clk, id_router_032:clk, id_router_033:clk, id_router_034:clk, id_router_035:clk, id_router_036:clk, id_router_037:clk, id_router_038:clk, id_router_039:clk, id_router_040:clk, id_router_041:clk, id_router_042:clk, id_router_043:clk, id_router_044:clk, id_router_045:clk, id_router_046:clk, id_router_047:clk, id_router_048:clk, id_router_049:clk, id_router_050:clk, id_router_051:clk, id_router_052:clk, id_router_053:clk, id_router_054:clk, id_router_055:clk, id_router_056:clk, id_router_057:clk, irq_mapper:clk, irq_synchronizer:receiver_clk, irq_synchronizer:sender_clk, limiter:clk, qsys_test_LEDState_0:csi_MCLK_clk, qsys_test_LEDState_1:csi_MCLK_clk, qsys_test_LEDState_2:csi_MCLK_clk, qsys_test_LEDState_3:csi_MCLK_clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_demux_019:clk, rsp_xbar_demux_020:clk, rsp_xbar_demux_021:clk, rsp_xbar_demux_022:clk, rsp_xbar_demux_023:clk, rsp_xbar_demux_024:clk, rsp_xbar_demux_025:clk, rsp_xbar_demux_026:clk, rsp_xbar_demux_027:clk, rsp_xbar_demux_028:clk, rsp_xbar_demux_029:clk, rsp_xbar_demux_030:clk, rsp_xbar_demux_031:clk, rsp_xbar_demux_032:clk, rsp_xbar_demux_033:clk, rsp_xbar_demux_034:clk, rsp_xbar_demux_035:clk, rsp_xbar_demux_036:clk, rsp_xbar_demux_037:clk, rsp_xbar_demux_038:clk, rsp_xbar_demux_039:clk, rsp_xbar_demux_040:clk, rsp_xbar_demux_041:clk, rsp_xbar_demux_042:clk, rsp_xbar_demux_043:clk, rsp_xbar_demux_044:clk, rsp_xbar_demux_045:clk, rsp_xbar_demux_046:clk, rsp_xbar_demux_047:clk, rsp_xbar_demux_048:clk, rsp_xbar_demux_049:clk, rsp_xbar_demux_050:clk, rsp_xbar_demux_051:clk, rsp_xbar_demux_052:clk, rsp_xbar_demux_053:clk, rsp_xbar_demux_054:clk, rsp_xbar_demux_055:clk, rsp_xbar_demux_056:clk, rsp_xbar_demux_057:clk, rsp_xbar_mux:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk, width_adapter_008:clk, width_adapter_009:clk, width_adapter_010:clk, width_adapter_011:clk, width_adapter_012:clk, width_adapter_013:clk, width_adapter_014:clk, width_adapter_015:clk, width_adapter_016:clk, width_adapter_017:clk, width_adapter_018:clk, width_adapter_019:clk, width_adapter_020:clk, width_adapter_021:clk, width_adapter_022:clk, width_adapter_023:clk, width_adapter_024:clk, width_adapter_025:clk, width_adapter_026:clk, width_adapter_027:clk, width_adapter_028:clk, width_adapter_029:clk, width_adapter_030:clk, width_adapter_031:clk, width_adapter_032:clk, width_adapter_033:clk, width_adapter_034:clk, width_adapter_035:clk, width_adapter_036:clk, width_adapter_037:clk, width_adapter_038:clk, width_adapter_039:clk, width_adapter_040:clk, width_adapter_041:clk, width_adapter_042:clk, width_adapter_043:clk, width_adapter_044:clk, width_adapter_045:clk, width_adapter_046:clk, width_adapter_047:clk, width_adapter_048:clk, width_adapter_049:clk, width_adapter_050:clk, width_adapter_051:clk, width_adapter_052:clk, width_adapter_053:clk, width_adapter_054:clk, width_adapter_055:clk, width_adapter_056:clk, width_adapter_057:clk, width_adapter_058:clk, width_adapter_059:clk, width_adapter_060:clk, width_adapter_061:clk, width_adapter_062:clk, width_adapter_063:clk, width_adapter_064:clk, width_adapter_065:clk, width_adapter_066:clk, width_adapter_067:clk, width_adapter_068:clk, width_adapter_069:clk, width_adapter_070:clk, width_adapter_071:clk, width_adapter_072:clk, width_adapter_073:clk, width_adapter_074:clk, width_adapter_075:clk, width_adapter_076:clk, width_adapter_077:clk, width_adapter_078:clk, width_adapter_079:clk, width_adapter_080:clk, width_adapter_081:clk, width_adapter_082:clk, width_adapter_083:clk, width_adapter_084:clk, width_adapter_085:clk, width_adapter_086:clk, width_adapter_087:clk, width_adapter_088:clk, width_adapter_089:clk, width_adapter_090:clk, width_adapter_091:clk, width_adapter_092:clk, width_adapter_093:clk, width_adapter_094:clk, width_adapter_095:clk, width_adapter_096:clk, width_adapter_097:clk, width_adapter_098:clk, width_adapter_099:clk, width_adapter_100:clk, width_adapter_101:clk, width_adapter_102:clk, width_adapter_103:clk]
	wire         qsys_test_ledstate_0_leds_valid;                                                         // qsys_test_LEDState_0:aso_LEDS_valid -> FuncLED_0:asi_LEDS_valid
	wire  [23:0] qsys_test_ledstate_0_leds_data;                                                          // qsys_test_LEDState_0:aso_LEDS_data -> FuncLED_0:asi_LEDS_data
	wire         qsys_test_ledstate_0_leds_ready;                                                         // FuncLED_0:asi_LEDS_ready -> qsys_test_LEDState_0:aso_LEDS_ready
	wire         qsys_test_ledstate_1_leds_valid;                                                         // qsys_test_LEDState_1:aso_LEDS_valid -> FuncLED_1:asi_LEDS_valid
	wire  [23:0] qsys_test_ledstate_1_leds_data;                                                          // qsys_test_LEDState_1:aso_LEDS_data -> FuncLED_1:asi_LEDS_data
	wire         qsys_test_ledstate_1_leds_ready;                                                         // FuncLED_1:asi_LEDS_ready -> qsys_test_LEDState_1:aso_LEDS_ready
	wire         qsys_test_ledstate_2_leds_valid;                                                         // qsys_test_LEDState_2:aso_LEDS_valid -> FuncLED_2:asi_LEDS_valid
	wire  [23:0] qsys_test_ledstate_2_leds_data;                                                          // qsys_test_LEDState_2:aso_LEDS_data -> FuncLED_2:asi_LEDS_data
	wire         qsys_test_ledstate_2_leds_ready;                                                         // FuncLED_2:asi_LEDS_ready -> qsys_test_LEDState_2:aso_LEDS_ready
	wire         qsys_test_ledstate_3_leds_valid;                                                         // qsys_test_LEDState_3:aso_LEDS_valid -> FuncLED_3:asi_LEDS_valid
	wire  [23:0] qsys_test_ledstate_3_leds_data;                                                          // qsys_test_LEDState_3:aso_LEDS_data -> FuncLED_3:asi_LEDS_data
	wire         qsys_test_ledstate_3_leds_ready;                                                         // FuncLED_3:asi_LEDS_ready -> qsys_test_LEDState_3:aso_LEDS_ready
	wire         sam9_m1_waitrequest;                                                                     // SAM9_M1_translator:av_waitrequest -> SAM9:avm_M1_waitrequest
	wire  [31:0] sam9_m1_address;                                                                         // SAM9:avm_M1_address -> SAM9_M1_translator:av_address
	wire  [31:0] sam9_m1_writedata;                                                                       // SAM9:avm_M1_writedata -> SAM9_M1_translator:av_writedata
	wire         sam9_m1_write;                                                                           // SAM9:avm_M1_write -> SAM9_M1_translator:av_write
	wire         sam9_m1_read;                                                                            // SAM9:avm_M1_read -> SAM9_M1_translator:av_read
	wire  [31:0] sam9_m1_readdata;                                                                        // SAM9_M1_translator:av_readdata -> SAM9:avm_M1_readdata
	wire         sam9_m1_begintransfer;                                                                   // SAM9:avm_M1_begintransfer -> SAM9_M1_translator:av_begintransfer
	wire         sam9_m1_readdatavalid;                                                                   // SAM9_M1_translator:av_readdatavalid -> SAM9:avm_M1_readdatavalid
	wire   [3:0] sam9_m1_byteenable;                                                                      // SAM9:avm_M1_byteenable -> SAM9_M1_translator:av_byteenable
	wire         sysid_sysid_translator_avalon_anti_slave_0_waitrequest;                                  // SysID:avs_SysID_waitrequest -> SysID_SysID_translator:av_waitrequest
	wire         sysid_sysid_translator_avalon_anti_slave_0_read;                                         // SysID_SysID_translator:av_read -> SysID:avs_SysID_read
	wire  [31:0] sysid_sysid_translator_avalon_anti_slave_0_readdata;                                     // SysID:avs_SysID_readdata -> SysID_SysID_translator:av_readdata
	wire         funcled_0_ledd_translator_avalon_anti_slave_0_waitrequest;                               // FuncLED_0:avs_LEDD_waitrequest -> FuncLED_0_LEDD_translator:av_waitrequest
	wire  [31:0] funcled_0_ledd_translator_avalon_anti_slave_0_writedata;                                 // FuncLED_0_LEDD_translator:av_writedata -> FuncLED_0:avs_LEDD_writedata
	wire         funcled_0_ledd_translator_avalon_anti_slave_0_write;                                     // FuncLED_0_LEDD_translator:av_write -> FuncLED_0:avs_LEDD_write
	wire         funcled_0_ledd_translator_avalon_anti_slave_0_read;                                      // FuncLED_0_LEDD_translator:av_read -> FuncLED_0:avs_LEDD_read
	wire  [31:0] funcled_0_ledd_translator_avalon_anti_slave_0_readdata;                                  // FuncLED_0:avs_LEDD_readdata -> FuncLED_0_LEDD_translator:av_readdata
	wire   [3:0] funcled_0_ledd_translator_avalon_anti_slave_0_byteenable;                                // FuncLED_0_LEDD_translator:av_byteenable -> FuncLED_0:avs_LEDD_byteenable
	wire         funcled_1_ledd_translator_avalon_anti_slave_0_waitrequest;                               // FuncLED_1:avs_LEDD_waitrequest -> FuncLED_1_LEDD_translator:av_waitrequest
	wire  [31:0] funcled_1_ledd_translator_avalon_anti_slave_0_writedata;                                 // FuncLED_1_LEDD_translator:av_writedata -> FuncLED_1:avs_LEDD_writedata
	wire         funcled_1_ledd_translator_avalon_anti_slave_0_write;                                     // FuncLED_1_LEDD_translator:av_write -> FuncLED_1:avs_LEDD_write
	wire         funcled_1_ledd_translator_avalon_anti_slave_0_read;                                      // FuncLED_1_LEDD_translator:av_read -> FuncLED_1:avs_LEDD_read
	wire  [31:0] funcled_1_ledd_translator_avalon_anti_slave_0_readdata;                                  // FuncLED_1:avs_LEDD_readdata -> FuncLED_1_LEDD_translator:av_readdata
	wire   [3:0] funcled_1_ledd_translator_avalon_anti_slave_0_byteenable;                                // FuncLED_1_LEDD_translator:av_byteenable -> FuncLED_1:avs_LEDD_byteenable
	wire         funcled_2_ledd_translator_avalon_anti_slave_0_waitrequest;                               // FuncLED_2:avs_LEDD_waitrequest -> FuncLED_2_LEDD_translator:av_waitrequest
	wire  [31:0] funcled_2_ledd_translator_avalon_anti_slave_0_writedata;                                 // FuncLED_2_LEDD_translator:av_writedata -> FuncLED_2:avs_LEDD_writedata
	wire         funcled_2_ledd_translator_avalon_anti_slave_0_write;                                     // FuncLED_2_LEDD_translator:av_write -> FuncLED_2:avs_LEDD_write
	wire         funcled_2_ledd_translator_avalon_anti_slave_0_read;                                      // FuncLED_2_LEDD_translator:av_read -> FuncLED_2:avs_LEDD_read
	wire  [31:0] funcled_2_ledd_translator_avalon_anti_slave_0_readdata;                                  // FuncLED_2:avs_LEDD_readdata -> FuncLED_2_LEDD_translator:av_readdata
	wire   [3:0] funcled_2_ledd_translator_avalon_anti_slave_0_byteenable;                                // FuncLED_2_LEDD_translator:av_byteenable -> FuncLED_2:avs_LEDD_byteenable
	wire         funcled_3_ledd_translator_avalon_anti_slave_0_waitrequest;                               // FuncLED_3:avs_LEDD_waitrequest -> FuncLED_3_LEDD_translator:av_waitrequest
	wire  [31:0] funcled_3_ledd_translator_avalon_anti_slave_0_writedata;                                 // FuncLED_3_LEDD_translator:av_writedata -> FuncLED_3:avs_LEDD_writedata
	wire         funcled_3_ledd_translator_avalon_anti_slave_0_write;                                     // FuncLED_3_LEDD_translator:av_write -> FuncLED_3:avs_LEDD_write
	wire         funcled_3_ledd_translator_avalon_anti_slave_0_read;                                      // FuncLED_3_LEDD_translator:av_read -> FuncLED_3:avs_LEDD_read
	wire  [31:0] funcled_3_ledd_translator_avalon_anti_slave_0_readdata;                                  // FuncLED_3:avs_LEDD_readdata -> FuncLED_3_LEDD_translator:av_readdata
	wire   [3:0] funcled_3_ledd_translator_avalon_anti_slave_0_byteenable;                                // FuncLED_3_LEDD_translator:av_byteenable -> FuncLED_3:avs_LEDD_byteenable
	wire         shield_admin_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shield_Admin:avs_Ctrl_waitrequest -> Shield_Admin_Ctrl_translator:av_waitrequest
	wire  [31:0] shield_admin_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shield_Admin_Ctrl_translator:av_writedata -> Shield_Admin:avs_Ctrl_writedata
	wire         shield_admin_ctrl_translator_avalon_anti_slave_0_write;                                  // Shield_Admin_Ctrl_translator:av_write -> Shield_Admin:avs_Ctrl_write
	wire         shield_admin_ctrl_translator_avalon_anti_slave_0_read;                                   // Shield_Admin_Ctrl_translator:av_read -> Shield_Admin:avs_Ctrl_read
	wire  [31:0] shield_admin_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shield_Admin:avs_Ctrl_readdata -> Shield_Admin_Ctrl_translator:av_readdata
	wire   [3:0] shield_admin_ctrl_translator_avalon_anti_slave_0_byteenable;                             // Shield_Admin_Ctrl_translator:av_byteenable -> Shield_Admin:avs_Ctrl_byteenable
	wire         shiled_io_a0_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_A0:avs_ctrl_waitrequest -> Shiled_IO_A0_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a0_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_A0_ctrl_translator:av_writedata -> Shiled_IO_A0:avs_ctrl_writedata
	wire         shiled_io_a0_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_A0_ctrl_translator:av_write -> Shiled_IO_A0:avs_ctrl_write
	wire         shiled_io_a0_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_A0_ctrl_translator:av_read -> Shiled_IO_A0:avs_ctrl_read
	wire   [7:0] shiled_io_a0_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_A0:avs_ctrl_readdata -> Shiled_IO_A0_ctrl_translator:av_readdata
	wire         shiled_io_a1_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_A1:avs_ctrl_waitrequest -> Shiled_IO_A1_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a1_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_A1_ctrl_translator:av_writedata -> Shiled_IO_A1:avs_ctrl_writedata
	wire         shiled_io_a1_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_A1_ctrl_translator:av_write -> Shiled_IO_A1:avs_ctrl_write
	wire         shiled_io_a1_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_A1_ctrl_translator:av_read -> Shiled_IO_A1:avs_ctrl_read
	wire   [7:0] shiled_io_a1_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_A1:avs_ctrl_readdata -> Shiled_IO_A1_ctrl_translator:av_readdata
	wire         shiled_io_a2_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_A2:avs_ctrl_waitrequest -> Shiled_IO_A2_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a2_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_A2_ctrl_translator:av_writedata -> Shiled_IO_A2:avs_ctrl_writedata
	wire         shiled_io_a2_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_A2_ctrl_translator:av_write -> Shiled_IO_A2:avs_ctrl_write
	wire         shiled_io_a2_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_A2_ctrl_translator:av_read -> Shiled_IO_A2:avs_ctrl_read
	wire   [7:0] shiled_io_a2_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_A2:avs_ctrl_readdata -> Shiled_IO_A2_ctrl_translator:av_readdata
	wire         shiled_io_a3_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_A3:avs_ctrl_waitrequest -> Shiled_IO_A3_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a3_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_A3_ctrl_translator:av_writedata -> Shiled_IO_A3:avs_ctrl_writedata
	wire         shiled_io_a3_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_A3_ctrl_translator:av_write -> Shiled_IO_A3:avs_ctrl_write
	wire         shiled_io_a3_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_A3_ctrl_translator:av_read -> Shiled_IO_A3:avs_ctrl_read
	wire   [7:0] shiled_io_a3_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_A3:avs_ctrl_readdata -> Shiled_IO_A3_ctrl_translator:av_readdata
	wire         shiled_io_a4_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_A4:avs_ctrl_waitrequest -> Shiled_IO_A4_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a4_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_A4_ctrl_translator:av_writedata -> Shiled_IO_A4:avs_ctrl_writedata
	wire         shiled_io_a4_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_A4_ctrl_translator:av_write -> Shiled_IO_A4:avs_ctrl_write
	wire         shiled_io_a4_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_A4_ctrl_translator:av_read -> Shiled_IO_A4:avs_ctrl_read
	wire   [7:0] shiled_io_a4_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_A4:avs_ctrl_readdata -> Shiled_IO_A4_ctrl_translator:av_readdata
	wire         shiled_io_a5_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_A5:avs_ctrl_waitrequest -> Shiled_IO_A5_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a5_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_A5_ctrl_translator:av_writedata -> Shiled_IO_A5:avs_ctrl_writedata
	wire         shiled_io_a5_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_A5_ctrl_translator:av_write -> Shiled_IO_A5:avs_ctrl_write
	wire         shiled_io_a5_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_A5_ctrl_translator:av_read -> Shiled_IO_A5:avs_ctrl_read
	wire   [7:0] shiled_io_a5_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_A5:avs_ctrl_readdata -> Shiled_IO_A5_ctrl_translator:av_readdata
	wire         shiled_io_a6_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_A6:avs_ctrl_waitrequest -> Shiled_IO_A6_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a6_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_A6_ctrl_translator:av_writedata -> Shiled_IO_A6:avs_ctrl_writedata
	wire         shiled_io_a6_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_A6_ctrl_translator:av_write -> Shiled_IO_A6:avs_ctrl_write
	wire         shiled_io_a6_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_A6_ctrl_translator:av_read -> Shiled_IO_A6:avs_ctrl_read
	wire   [7:0] shiled_io_a6_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_A6:avs_ctrl_readdata -> Shiled_IO_A6_ctrl_translator:av_readdata
	wire         shiled_io_a7_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_A7:avs_ctrl_waitrequest -> Shiled_IO_A7_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a7_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_A7_ctrl_translator:av_writedata -> Shiled_IO_A7:avs_ctrl_writedata
	wire         shiled_io_a7_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_A7_ctrl_translator:av_write -> Shiled_IO_A7:avs_ctrl_write
	wire         shiled_io_a7_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_A7_ctrl_translator:av_read -> Shiled_IO_A7:avs_ctrl_read
	wire   [7:0] shiled_io_a7_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_A7:avs_ctrl_readdata -> Shiled_IO_A7_ctrl_translator:av_readdata
	wire         shiled_io_a8_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_A8:avs_ctrl_waitrequest -> Shiled_IO_A8_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a8_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_A8_ctrl_translator:av_writedata -> Shiled_IO_A8:avs_ctrl_writedata
	wire         shiled_io_a8_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_A8_ctrl_translator:av_write -> Shiled_IO_A8:avs_ctrl_write
	wire         shiled_io_a8_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_A8_ctrl_translator:av_read -> Shiled_IO_A8:avs_ctrl_read
	wire   [7:0] shiled_io_a8_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_A8:avs_ctrl_readdata -> Shiled_IO_A8_ctrl_translator:av_readdata
	wire         shiled_io_a9_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_A9:avs_ctrl_waitrequest -> Shiled_IO_A9_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a9_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_A9_ctrl_translator:av_writedata -> Shiled_IO_A9:avs_ctrl_writedata
	wire         shiled_io_a9_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_A9_ctrl_translator:av_write -> Shiled_IO_A9:avs_ctrl_write
	wire         shiled_io_a9_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_A9_ctrl_translator:av_read -> Shiled_IO_A9:avs_ctrl_read
	wire   [7:0] shiled_io_a9_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_A9:avs_ctrl_readdata -> Shiled_IO_A9_ctrl_translator:av_readdata
	wire         shiled_io_a10_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A10:avs_ctrl_waitrequest -> Shiled_IO_A10_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a10_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A10_ctrl_translator:av_writedata -> Shiled_IO_A10:avs_ctrl_writedata
	wire         shiled_io_a10_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A10_ctrl_translator:av_write -> Shiled_IO_A10:avs_ctrl_write
	wire         shiled_io_a10_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A10_ctrl_translator:av_read -> Shiled_IO_A10:avs_ctrl_read
	wire   [7:0] shiled_io_a10_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A10:avs_ctrl_readdata -> Shiled_IO_A10_ctrl_translator:av_readdata
	wire         shiled_io_a11_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A11:avs_ctrl_waitrequest -> Shiled_IO_A11_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a11_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A11_ctrl_translator:av_writedata -> Shiled_IO_A11:avs_ctrl_writedata
	wire         shiled_io_a11_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A11_ctrl_translator:av_write -> Shiled_IO_A11:avs_ctrl_write
	wire         shiled_io_a11_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A11_ctrl_translator:av_read -> Shiled_IO_A11:avs_ctrl_read
	wire   [7:0] shiled_io_a11_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A11:avs_ctrl_readdata -> Shiled_IO_A11_ctrl_translator:av_readdata
	wire         shiled_io_a13_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A13:avs_ctrl_waitrequest -> Shiled_IO_A13_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a13_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A13_ctrl_translator:av_writedata -> Shiled_IO_A13:avs_ctrl_writedata
	wire         shiled_io_a13_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A13_ctrl_translator:av_write -> Shiled_IO_A13:avs_ctrl_write
	wire         shiled_io_a13_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A13_ctrl_translator:av_read -> Shiled_IO_A13:avs_ctrl_read
	wire   [7:0] shiled_io_a13_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A13:avs_ctrl_readdata -> Shiled_IO_A13_ctrl_translator:av_readdata
	wire         shiled_io_a12_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A12:avs_ctrl_waitrequest -> Shiled_IO_A12_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a12_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A12_ctrl_translator:av_writedata -> Shiled_IO_A12:avs_ctrl_writedata
	wire         shiled_io_a12_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A12_ctrl_translator:av_write -> Shiled_IO_A12:avs_ctrl_write
	wire         shiled_io_a12_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A12_ctrl_translator:av_read -> Shiled_IO_A12:avs_ctrl_read
	wire   [7:0] shiled_io_a12_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A12:avs_ctrl_readdata -> Shiled_IO_A12_ctrl_translator:av_readdata
	wire         shiled_io_a14_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A14:avs_ctrl_waitrequest -> Shiled_IO_A14_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a14_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A14_ctrl_translator:av_writedata -> Shiled_IO_A14:avs_ctrl_writedata
	wire         shiled_io_a14_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A14_ctrl_translator:av_write -> Shiled_IO_A14:avs_ctrl_write
	wire         shiled_io_a14_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A14_ctrl_translator:av_read -> Shiled_IO_A14:avs_ctrl_read
	wire   [7:0] shiled_io_a14_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A14:avs_ctrl_readdata -> Shiled_IO_A14_ctrl_translator:av_readdata
	wire         shiled_io_a15_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A15:avs_ctrl_waitrequest -> Shiled_IO_A15_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a15_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A15_ctrl_translator:av_writedata -> Shiled_IO_A15:avs_ctrl_writedata
	wire         shiled_io_a15_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A15_ctrl_translator:av_write -> Shiled_IO_A15:avs_ctrl_write
	wire         shiled_io_a15_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A15_ctrl_translator:av_read -> Shiled_IO_A15:avs_ctrl_read
	wire   [7:0] shiled_io_a15_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A15:avs_ctrl_readdata -> Shiled_IO_A15_ctrl_translator:av_readdata
	wire         shiled_io_a17_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A17:avs_ctrl_waitrequest -> Shiled_IO_A17_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a17_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A17_ctrl_translator:av_writedata -> Shiled_IO_A17:avs_ctrl_writedata
	wire         shiled_io_a17_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A17_ctrl_translator:av_write -> Shiled_IO_A17:avs_ctrl_write
	wire         shiled_io_a17_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A17_ctrl_translator:av_read -> Shiled_IO_A17:avs_ctrl_read
	wire   [7:0] shiled_io_a17_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A17:avs_ctrl_readdata -> Shiled_IO_A17_ctrl_translator:av_readdata
	wire         shiled_io_a16_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A16:avs_ctrl_waitrequest -> Shiled_IO_A16_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a16_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A16_ctrl_translator:av_writedata -> Shiled_IO_A16:avs_ctrl_writedata
	wire         shiled_io_a16_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A16_ctrl_translator:av_write -> Shiled_IO_A16:avs_ctrl_write
	wire         shiled_io_a16_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A16_ctrl_translator:av_read -> Shiled_IO_A16:avs_ctrl_read
	wire   [7:0] shiled_io_a16_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A16:avs_ctrl_readdata -> Shiled_IO_A16_ctrl_translator:av_readdata
	wire         shiled_io_a18_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A18:avs_ctrl_waitrequest -> Shiled_IO_A18_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a18_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A18_ctrl_translator:av_writedata -> Shiled_IO_A18:avs_ctrl_writedata
	wire         shiled_io_a18_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A18_ctrl_translator:av_write -> Shiled_IO_A18:avs_ctrl_write
	wire         shiled_io_a18_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A18_ctrl_translator:av_read -> Shiled_IO_A18:avs_ctrl_read
	wire   [7:0] shiled_io_a18_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A18:avs_ctrl_readdata -> Shiled_IO_A18_ctrl_translator:av_readdata
	wire         shiled_io_a19_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A19:avs_ctrl_waitrequest -> Shiled_IO_A19_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a19_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A19_ctrl_translator:av_writedata -> Shiled_IO_A19:avs_ctrl_writedata
	wire         shiled_io_a19_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A19_ctrl_translator:av_write -> Shiled_IO_A19:avs_ctrl_write
	wire         shiled_io_a19_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A19_ctrl_translator:av_read -> Shiled_IO_A19:avs_ctrl_read
	wire   [7:0] shiled_io_a19_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A19:avs_ctrl_readdata -> Shiled_IO_A19_ctrl_translator:av_readdata
	wire         shiled_io_a20_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A20:avs_ctrl_waitrequest -> Shiled_IO_A20_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a20_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A20_ctrl_translator:av_writedata -> Shiled_IO_A20:avs_ctrl_writedata
	wire         shiled_io_a20_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A20_ctrl_translator:av_write -> Shiled_IO_A20:avs_ctrl_write
	wire         shiled_io_a20_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A20_ctrl_translator:av_read -> Shiled_IO_A20:avs_ctrl_read
	wire   [7:0] shiled_io_a20_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A20:avs_ctrl_readdata -> Shiled_IO_A20_ctrl_translator:av_readdata
	wire         shiled_io_a21_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A21:avs_ctrl_waitrequest -> Shiled_IO_A21_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a21_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A21_ctrl_translator:av_writedata -> Shiled_IO_A21:avs_ctrl_writedata
	wire         shiled_io_a21_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A21_ctrl_translator:av_write -> Shiled_IO_A21:avs_ctrl_write
	wire         shiled_io_a21_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A21_ctrl_translator:av_read -> Shiled_IO_A21:avs_ctrl_read
	wire   [7:0] shiled_io_a21_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A21:avs_ctrl_readdata -> Shiled_IO_A21_ctrl_translator:av_readdata
	wire         shiled_io_a22_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A22:avs_ctrl_waitrequest -> Shiled_IO_A22_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a22_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A22_ctrl_translator:av_writedata -> Shiled_IO_A22:avs_ctrl_writedata
	wire         shiled_io_a22_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A22_ctrl_translator:av_write -> Shiled_IO_A22:avs_ctrl_write
	wire         shiled_io_a22_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A22_ctrl_translator:av_read -> Shiled_IO_A22:avs_ctrl_read
	wire   [7:0] shiled_io_a22_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A22:avs_ctrl_readdata -> Shiled_IO_A22_ctrl_translator:av_readdata
	wire         shiled_io_a23_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A23:avs_ctrl_waitrequest -> Shiled_IO_A23_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a23_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A23_ctrl_translator:av_writedata -> Shiled_IO_A23:avs_ctrl_writedata
	wire         shiled_io_a23_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A23_ctrl_translator:av_write -> Shiled_IO_A23:avs_ctrl_write
	wire         shiled_io_a23_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A23_ctrl_translator:av_read -> Shiled_IO_A23:avs_ctrl_read
	wire   [7:0] shiled_io_a23_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A23:avs_ctrl_readdata -> Shiled_IO_A23_ctrl_translator:av_readdata
	wire         shiled_io_a24_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A24:avs_ctrl_waitrequest -> Shiled_IO_A24_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a24_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A24_ctrl_translator:av_writedata -> Shiled_IO_A24:avs_ctrl_writedata
	wire         shiled_io_a24_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A24_ctrl_translator:av_write -> Shiled_IO_A24:avs_ctrl_write
	wire         shiled_io_a24_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A24_ctrl_translator:av_read -> Shiled_IO_A24:avs_ctrl_read
	wire   [7:0] shiled_io_a24_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A24:avs_ctrl_readdata -> Shiled_IO_A24_ctrl_translator:av_readdata
	wire         shiled_io_a25_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_A25:avs_ctrl_waitrequest -> Shiled_IO_A25_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_a25_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_A25_ctrl_translator:av_writedata -> Shiled_IO_A25:avs_ctrl_writedata
	wire         shiled_io_a25_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_A25_ctrl_translator:av_write -> Shiled_IO_A25:avs_ctrl_write
	wire         shiled_io_a25_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_A25_ctrl_translator:av_read -> Shiled_IO_A25:avs_ctrl_read
	wire   [7:0] shiled_io_a25_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_A25:avs_ctrl_readdata -> Shiled_IO_A25_ctrl_translator:av_readdata
	wire         shiled_io_b0_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_B0:avs_ctrl_waitrequest -> Shiled_IO_B0_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b0_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_B0_ctrl_translator:av_writedata -> Shiled_IO_B0:avs_ctrl_writedata
	wire         shiled_io_b0_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_B0_ctrl_translator:av_write -> Shiled_IO_B0:avs_ctrl_write
	wire         shiled_io_b0_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_B0_ctrl_translator:av_read -> Shiled_IO_B0:avs_ctrl_read
	wire   [7:0] shiled_io_b0_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_B0:avs_ctrl_readdata -> Shiled_IO_B0_ctrl_translator:av_readdata
	wire         shiled_io_b1_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_B1:avs_ctrl_waitrequest -> Shiled_IO_B1_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b1_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_B1_ctrl_translator:av_writedata -> Shiled_IO_B1:avs_ctrl_writedata
	wire         shiled_io_b1_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_B1_ctrl_translator:av_write -> Shiled_IO_B1:avs_ctrl_write
	wire         shiled_io_b1_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_B1_ctrl_translator:av_read -> Shiled_IO_B1:avs_ctrl_read
	wire   [7:0] shiled_io_b1_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_B1:avs_ctrl_readdata -> Shiled_IO_B1_ctrl_translator:av_readdata
	wire         shiled_io_b2_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_B2:avs_ctrl_waitrequest -> Shiled_IO_B2_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b2_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_B2_ctrl_translator:av_writedata -> Shiled_IO_B2:avs_ctrl_writedata
	wire         shiled_io_b2_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_B2_ctrl_translator:av_write -> Shiled_IO_B2:avs_ctrl_write
	wire         shiled_io_b2_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_B2_ctrl_translator:av_read -> Shiled_IO_B2:avs_ctrl_read
	wire   [7:0] shiled_io_b2_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_B2:avs_ctrl_readdata -> Shiled_IO_B2_ctrl_translator:av_readdata
	wire         shiled_io_b3_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_B3:avs_ctrl_waitrequest -> Shiled_IO_B3_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b3_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_B3_ctrl_translator:av_writedata -> Shiled_IO_B3:avs_ctrl_writedata
	wire         shiled_io_b3_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_B3_ctrl_translator:av_write -> Shiled_IO_B3:avs_ctrl_write
	wire         shiled_io_b3_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_B3_ctrl_translator:av_read -> Shiled_IO_B3:avs_ctrl_read
	wire   [7:0] shiled_io_b3_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_B3:avs_ctrl_readdata -> Shiled_IO_B3_ctrl_translator:av_readdata
	wire         shiled_io_b4_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_B4:avs_ctrl_waitrequest -> Shiled_IO_B4_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b4_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_B4_ctrl_translator:av_writedata -> Shiled_IO_B4:avs_ctrl_writedata
	wire         shiled_io_b4_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_B4_ctrl_translator:av_write -> Shiled_IO_B4:avs_ctrl_write
	wire         shiled_io_b4_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_B4_ctrl_translator:av_read -> Shiled_IO_B4:avs_ctrl_read
	wire   [7:0] shiled_io_b4_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_B4:avs_ctrl_readdata -> Shiled_IO_B4_ctrl_translator:av_readdata
	wire         shiled_io_b6_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_B6:avs_ctrl_waitrequest -> Shiled_IO_B6_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b6_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_B6_ctrl_translator:av_writedata -> Shiled_IO_B6:avs_ctrl_writedata
	wire         shiled_io_b6_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_B6_ctrl_translator:av_write -> Shiled_IO_B6:avs_ctrl_write
	wire         shiled_io_b6_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_B6_ctrl_translator:av_read -> Shiled_IO_B6:avs_ctrl_read
	wire   [7:0] shiled_io_b6_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_B6:avs_ctrl_readdata -> Shiled_IO_B6_ctrl_translator:av_readdata
	wire         shiled_io_b5_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_B5:avs_ctrl_waitrequest -> Shiled_IO_B5_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b5_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_B5_ctrl_translator:av_writedata -> Shiled_IO_B5:avs_ctrl_writedata
	wire         shiled_io_b5_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_B5_ctrl_translator:av_write -> Shiled_IO_B5:avs_ctrl_write
	wire         shiled_io_b5_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_B5_ctrl_translator:av_read -> Shiled_IO_B5:avs_ctrl_read
	wire   [7:0] shiled_io_b5_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_B5:avs_ctrl_readdata -> Shiled_IO_B5_ctrl_translator:av_readdata
	wire         shiled_io_b7_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_B7:avs_ctrl_waitrequest -> Shiled_IO_B7_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b7_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_B7_ctrl_translator:av_writedata -> Shiled_IO_B7:avs_ctrl_writedata
	wire         shiled_io_b7_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_B7_ctrl_translator:av_write -> Shiled_IO_B7:avs_ctrl_write
	wire         shiled_io_b7_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_B7_ctrl_translator:av_read -> Shiled_IO_B7:avs_ctrl_read
	wire   [7:0] shiled_io_b7_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_B7:avs_ctrl_readdata -> Shiled_IO_B7_ctrl_translator:av_readdata
	wire         shiled_io_b8_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_B8:avs_ctrl_waitrequest -> Shiled_IO_B8_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b8_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_B8_ctrl_translator:av_writedata -> Shiled_IO_B8:avs_ctrl_writedata
	wire         shiled_io_b8_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_B8_ctrl_translator:av_write -> Shiled_IO_B8:avs_ctrl_write
	wire         shiled_io_b8_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_B8_ctrl_translator:av_read -> Shiled_IO_B8:avs_ctrl_read
	wire   [7:0] shiled_io_b8_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_B8:avs_ctrl_readdata -> Shiled_IO_B8_ctrl_translator:av_readdata
	wire         shiled_io_b9_ctrl_translator_avalon_anti_slave_0_waitrequest;                            // Shiled_IO_B9:avs_ctrl_waitrequest -> Shiled_IO_B9_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b9_ctrl_translator_avalon_anti_slave_0_writedata;                              // Shiled_IO_B9_ctrl_translator:av_writedata -> Shiled_IO_B9:avs_ctrl_writedata
	wire         shiled_io_b9_ctrl_translator_avalon_anti_slave_0_write;                                  // Shiled_IO_B9_ctrl_translator:av_write -> Shiled_IO_B9:avs_ctrl_write
	wire         shiled_io_b9_ctrl_translator_avalon_anti_slave_0_read;                                   // Shiled_IO_B9_ctrl_translator:av_read -> Shiled_IO_B9:avs_ctrl_read
	wire   [7:0] shiled_io_b9_ctrl_translator_avalon_anti_slave_0_readdata;                               // Shiled_IO_B9:avs_ctrl_readdata -> Shiled_IO_B9_ctrl_translator:av_readdata
	wire         shiled_io_b10_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B10:avs_ctrl_waitrequest -> Shiled_IO_B10_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b10_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B10_ctrl_translator:av_writedata -> Shiled_IO_B10:avs_ctrl_writedata
	wire         shiled_io_b10_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B10_ctrl_translator:av_write -> Shiled_IO_B10:avs_ctrl_write
	wire         shiled_io_b10_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B10_ctrl_translator:av_read -> Shiled_IO_B10:avs_ctrl_read
	wire   [7:0] shiled_io_b10_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B10:avs_ctrl_readdata -> Shiled_IO_B10_ctrl_translator:av_readdata
	wire         shiled_io_b11_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B11:avs_ctrl_waitrequest -> Shiled_IO_B11_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b11_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B11_ctrl_translator:av_writedata -> Shiled_IO_B11:avs_ctrl_writedata
	wire         shiled_io_b11_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B11_ctrl_translator:av_write -> Shiled_IO_B11:avs_ctrl_write
	wire         shiled_io_b11_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B11_ctrl_translator:av_read -> Shiled_IO_B11:avs_ctrl_read
	wire   [7:0] shiled_io_b11_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B11:avs_ctrl_readdata -> Shiled_IO_B11_ctrl_translator:av_readdata
	wire         shiled_io_b12_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B12:avs_ctrl_waitrequest -> Shiled_IO_B12_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b12_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B12_ctrl_translator:av_writedata -> Shiled_IO_B12:avs_ctrl_writedata
	wire         shiled_io_b12_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B12_ctrl_translator:av_write -> Shiled_IO_B12:avs_ctrl_write
	wire         shiled_io_b12_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B12_ctrl_translator:av_read -> Shiled_IO_B12:avs_ctrl_read
	wire   [7:0] shiled_io_b12_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B12:avs_ctrl_readdata -> Shiled_IO_B12_ctrl_translator:av_readdata
	wire         shiled_io_b13_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B13:avs_ctrl_waitrequest -> Shiled_IO_B13_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b13_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B13_ctrl_translator:av_writedata -> Shiled_IO_B13:avs_ctrl_writedata
	wire         shiled_io_b13_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B13_ctrl_translator:av_write -> Shiled_IO_B13:avs_ctrl_write
	wire         shiled_io_b13_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B13_ctrl_translator:av_read -> Shiled_IO_B13:avs_ctrl_read
	wire   [7:0] shiled_io_b13_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B13:avs_ctrl_readdata -> Shiled_IO_B13_ctrl_translator:av_readdata
	wire         shiled_io_b14_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B14:avs_ctrl_waitrequest -> Shiled_IO_B14_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b14_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B14_ctrl_translator:av_writedata -> Shiled_IO_B14:avs_ctrl_writedata
	wire         shiled_io_b14_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B14_ctrl_translator:av_write -> Shiled_IO_B14:avs_ctrl_write
	wire         shiled_io_b14_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B14_ctrl_translator:av_read -> Shiled_IO_B14:avs_ctrl_read
	wire   [7:0] shiled_io_b14_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B14:avs_ctrl_readdata -> Shiled_IO_B14_ctrl_translator:av_readdata
	wire         shiled_io_b15_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B15:avs_ctrl_waitrequest -> Shiled_IO_B15_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b15_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B15_ctrl_translator:av_writedata -> Shiled_IO_B15:avs_ctrl_writedata
	wire         shiled_io_b15_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B15_ctrl_translator:av_write -> Shiled_IO_B15:avs_ctrl_write
	wire         shiled_io_b15_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B15_ctrl_translator:av_read -> Shiled_IO_B15:avs_ctrl_read
	wire   [7:0] shiled_io_b15_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B15:avs_ctrl_readdata -> Shiled_IO_B15_ctrl_translator:av_readdata
	wire         shiled_io_b16_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B16:avs_ctrl_waitrequest -> Shiled_IO_B16_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b16_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B16_ctrl_translator:av_writedata -> Shiled_IO_B16:avs_ctrl_writedata
	wire         shiled_io_b16_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B16_ctrl_translator:av_write -> Shiled_IO_B16:avs_ctrl_write
	wire         shiled_io_b16_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B16_ctrl_translator:av_read -> Shiled_IO_B16:avs_ctrl_read
	wire   [7:0] shiled_io_b16_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B16:avs_ctrl_readdata -> Shiled_IO_B16_ctrl_translator:av_readdata
	wire         shiled_io_b17_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B17:avs_ctrl_waitrequest -> Shiled_IO_B17_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b17_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B17_ctrl_translator:av_writedata -> Shiled_IO_B17:avs_ctrl_writedata
	wire         shiled_io_b17_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B17_ctrl_translator:av_write -> Shiled_IO_B17:avs_ctrl_write
	wire         shiled_io_b17_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B17_ctrl_translator:av_read -> Shiled_IO_B17:avs_ctrl_read
	wire   [7:0] shiled_io_b17_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B17:avs_ctrl_readdata -> Shiled_IO_B17_ctrl_translator:av_readdata
	wire         shiled_io_b18_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B18:avs_ctrl_waitrequest -> Shiled_IO_B18_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b18_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B18_ctrl_translator:av_writedata -> Shiled_IO_B18:avs_ctrl_writedata
	wire         shiled_io_b18_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B18_ctrl_translator:av_write -> Shiled_IO_B18:avs_ctrl_write
	wire         shiled_io_b18_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B18_ctrl_translator:av_read -> Shiled_IO_B18:avs_ctrl_read
	wire   [7:0] shiled_io_b18_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B18:avs_ctrl_readdata -> Shiled_IO_B18_ctrl_translator:av_readdata
	wire         shiled_io_b19_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B19:avs_ctrl_waitrequest -> Shiled_IO_B19_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b19_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B19_ctrl_translator:av_writedata -> Shiled_IO_B19:avs_ctrl_writedata
	wire         shiled_io_b19_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B19_ctrl_translator:av_write -> Shiled_IO_B19:avs_ctrl_write
	wire         shiled_io_b19_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B19_ctrl_translator:av_read -> Shiled_IO_B19:avs_ctrl_read
	wire   [7:0] shiled_io_b19_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B19:avs_ctrl_readdata -> Shiled_IO_B19_ctrl_translator:av_readdata
	wire         shiled_io_b20_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B20:avs_ctrl_waitrequest -> Shiled_IO_B20_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b20_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B20_ctrl_translator:av_writedata -> Shiled_IO_B20:avs_ctrl_writedata
	wire         shiled_io_b20_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B20_ctrl_translator:av_write -> Shiled_IO_B20:avs_ctrl_write
	wire         shiled_io_b20_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B20_ctrl_translator:av_read -> Shiled_IO_B20:avs_ctrl_read
	wire   [7:0] shiled_io_b20_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B20:avs_ctrl_readdata -> Shiled_IO_B20_ctrl_translator:av_readdata
	wire         shiled_io_b21_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B21:avs_ctrl_waitrequest -> Shiled_IO_B21_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b21_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B21_ctrl_translator:av_writedata -> Shiled_IO_B21:avs_ctrl_writedata
	wire         shiled_io_b21_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B21_ctrl_translator:av_write -> Shiled_IO_B21:avs_ctrl_write
	wire         shiled_io_b21_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B21_ctrl_translator:av_read -> Shiled_IO_B21:avs_ctrl_read
	wire   [7:0] shiled_io_b21_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B21:avs_ctrl_readdata -> Shiled_IO_B21_ctrl_translator:av_readdata
	wire         shiled_io_b22_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B22:avs_ctrl_waitrequest -> Shiled_IO_B22_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b22_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B22_ctrl_translator:av_writedata -> Shiled_IO_B22:avs_ctrl_writedata
	wire         shiled_io_b22_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B22_ctrl_translator:av_write -> Shiled_IO_B22:avs_ctrl_write
	wire         shiled_io_b22_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B22_ctrl_translator:av_read -> Shiled_IO_B22:avs_ctrl_read
	wire   [7:0] shiled_io_b22_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B22:avs_ctrl_readdata -> Shiled_IO_B22_ctrl_translator:av_readdata
	wire         shiled_io_b23_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B23:avs_ctrl_waitrequest -> Shiled_IO_B23_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b23_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B23_ctrl_translator:av_writedata -> Shiled_IO_B23:avs_ctrl_writedata
	wire         shiled_io_b23_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B23_ctrl_translator:av_write -> Shiled_IO_B23:avs_ctrl_write
	wire         shiled_io_b23_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B23_ctrl_translator:av_read -> Shiled_IO_B23:avs_ctrl_read
	wire   [7:0] shiled_io_b23_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B23:avs_ctrl_readdata -> Shiled_IO_B23_ctrl_translator:av_readdata
	wire         shiled_io_b24_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B24:avs_ctrl_waitrequest -> Shiled_IO_B24_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b24_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B24_ctrl_translator:av_writedata -> Shiled_IO_B24:avs_ctrl_writedata
	wire         shiled_io_b24_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B24_ctrl_translator:av_write -> Shiled_IO_B24:avs_ctrl_write
	wire         shiled_io_b24_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B24_ctrl_translator:av_read -> Shiled_IO_B24:avs_ctrl_read
	wire   [7:0] shiled_io_b24_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B24:avs_ctrl_readdata -> Shiled_IO_B24_ctrl_translator:av_readdata
	wire         shiled_io_b25_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shiled_IO_B25:avs_ctrl_waitrequest -> Shiled_IO_B25_ctrl_translator:av_waitrequest
	wire   [7:0] shiled_io_b25_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shiled_IO_B25_ctrl_translator:av_writedata -> Shiled_IO_B25:avs_ctrl_writedata
	wire         shiled_io_b25_ctrl_translator_avalon_anti_slave_0_write;                                 // Shiled_IO_B25_ctrl_translator:av_write -> Shiled_IO_B25:avs_ctrl_write
	wire         shiled_io_b25_ctrl_translator_avalon_anti_slave_0_read;                                  // Shiled_IO_B25_ctrl_translator:av_read -> Shiled_IO_B25:avs_ctrl_read
	wire   [7:0] shiled_io_b25_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shiled_IO_B25:avs_ctrl_readdata -> Shiled_IO_B25_ctrl_translator:av_readdata
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_B0_ctrl_translator:uav_waitrequest -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B0_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B0_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B0_ctrl_translator:uav_address
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B0_ctrl_translator:uav_write
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B0_ctrl_translator:uav_lock
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B0_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_B0_ctrl_translator:uav_readdata -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_B0_ctrl_translator:uav_readdatavalid -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B0_ctrl_translator:uav_debugaccess
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B0_ctrl_translator:uav_byteenable
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_B2_ctrl_translator:uav_waitrequest -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B2_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B2_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B2_ctrl_translator:uav_address
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B2_ctrl_translator:uav_write
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B2_ctrl_translator:uav_lock
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B2_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_B2_ctrl_translator:uav_readdata -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_B2_ctrl_translator:uav_readdatavalid -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B2_ctrl_translator:uav_debugaccess
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B2_ctrl_translator:uav_byteenable
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A12_ctrl_translator:uav_waitrequest -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A12_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A12_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A12_ctrl_translator:uav_address
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A12_ctrl_translator:uav_write
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A12_ctrl_translator:uav_lock
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A12_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A12_ctrl_translator:uav_readdata -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A12_ctrl_translator:uav_readdatavalid -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A12_ctrl_translator:uav_debugaccess
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A12_ctrl_translator:uav_byteenable
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A11_ctrl_translator:uav_waitrequest -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A11_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A11_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A11_ctrl_translator:uav_address
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A11_ctrl_translator:uav_write
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A11_ctrl_translator:uav_lock
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A11_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A11_ctrl_translator:uav_readdata -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A11_ctrl_translator:uav_readdatavalid -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A11_ctrl_translator:uav_debugaccess
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A11_ctrl_translator:uav_byteenable
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_A1_ctrl_translator:uav_waitrequest -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A1_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A1_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A1_ctrl_translator:uav_address
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A1_ctrl_translator:uav_write
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A1_ctrl_translator:uav_lock
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A1_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_A1_ctrl_translator:uav_readdata -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_A1_ctrl_translator:uav_readdatavalid -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A1_ctrl_translator:uav_debugaccess
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A1_ctrl_translator:uav_byteenable
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_A0_ctrl_translator:uav_waitrequest -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A0_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A0_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A0_ctrl_translator:uav_address
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A0_ctrl_translator:uav_write
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A0_ctrl_translator:uav_lock
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A0_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_A0_ctrl_translator:uav_readdata -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_A0_ctrl_translator:uav_readdatavalid -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A0_ctrl_translator:uav_debugaccess
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A0_ctrl_translator:uav_byteenable
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B19_ctrl_translator:uav_waitrequest -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B19_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B19_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B19_ctrl_translator:uav_address
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B19_ctrl_translator:uav_write
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B19_ctrl_translator:uav_lock
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B19_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B19_ctrl_translator:uav_readdata -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B19_ctrl_translator:uav_readdatavalid -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B19_ctrl_translator:uav_debugaccess
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B19_ctrl_translator:uav_byteenable
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A10_ctrl_translator:uav_waitrequest -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A10_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A10_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A10_ctrl_translator:uav_address
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A10_ctrl_translator:uav_write
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A10_ctrl_translator:uav_lock
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A10_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A10_ctrl_translator:uav_readdata -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A10_ctrl_translator:uav_readdatavalid -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A10_ctrl_translator:uav_debugaccess
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A10_ctrl_translator:uav_byteenable
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A19_ctrl_translator:uav_waitrequest -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A19_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A19_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A19_ctrl_translator:uav_address
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A19_ctrl_translator:uav_write
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A19_ctrl_translator:uav_lock
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A19_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A19_ctrl_translator:uav_readdata -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A19_ctrl_translator:uav_readdatavalid -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A19_ctrl_translator:uav_debugaccess
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A19_ctrl_translator:uav_byteenable
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_B1_ctrl_translator:uav_waitrequest -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B1_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B1_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B1_ctrl_translator:uav_address
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B1_ctrl_translator:uav_write
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B1_ctrl_translator:uav_lock
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B1_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_B1_ctrl_translator:uav_readdata -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_B1_ctrl_translator:uav_readdatavalid -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B1_ctrl_translator:uav_debugaccess
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B1_ctrl_translator:uav_byteenable
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // FuncLED_0_LEDD_translator:uav_waitrequest -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> FuncLED_0_LEDD_translator:uav_burstcount
	wire  [31:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                   // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> FuncLED_0_LEDD_translator:uav_writedata
	wire  [31:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_address;                     // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> FuncLED_0_LEDD_translator:uav_address
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_write;                       // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> FuncLED_0_LEDD_translator:uav_write
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                        // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> FuncLED_0_LEDD_translator:uav_lock
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_read;                        // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> FuncLED_0_LEDD_translator:uav_read
	wire  [31:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                    // FuncLED_0_LEDD_translator:uav_readdata -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // FuncLED_0_LEDD_translator:uav_readdatavalid -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FuncLED_0_LEDD_translator:uav_debugaccess
	wire   [3:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> FuncLED_0_LEDD_translator:uav_byteenable
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;                // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                 // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;                // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_A6_ctrl_translator:uav_waitrequest -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A6_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A6_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A6_ctrl_translator:uav_address
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A6_ctrl_translator:uav_write
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A6_ctrl_translator:uav_lock
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A6_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_A6_ctrl_translator:uav_readdata -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_A6_ctrl_translator:uav_readdatavalid -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A6_ctrl_translator:uav_debugaccess
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A6_ctrl_translator:uav_byteenable
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_A4_ctrl_translator:uav_waitrequest -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A4_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A4_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A4_ctrl_translator:uav_address
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A4_ctrl_translator:uav_write
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A4_ctrl_translator:uav_lock
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A4_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_A4_ctrl_translator:uav_readdata -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_A4_ctrl_translator:uav_readdatavalid -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A4_ctrl_translator:uav_debugaccess
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A4_ctrl_translator:uav_byteenable
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A20_ctrl_translator:uav_waitrequest -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A20_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A20_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A20_ctrl_translator:uav_address
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A20_ctrl_translator:uav_write
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A20_ctrl_translator:uav_lock
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A20_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A20_ctrl_translator:uav_readdata -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A20_ctrl_translator:uav_readdatavalid -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A20_ctrl_translator:uav_debugaccess
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A20_ctrl_translator:uav_byteenable
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B11_ctrl_translator:uav_waitrequest -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B11_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B11_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B11_ctrl_translator:uav_address
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B11_ctrl_translator:uav_write
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B11_ctrl_translator:uav_lock
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B11_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B11_ctrl_translator:uav_readdata -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B11_ctrl_translator:uav_readdatavalid -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B11_ctrl_translator:uav_debugaccess
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B11_ctrl_translator:uav_byteenable
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A17_ctrl_translator:uav_waitrequest -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A17_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A17_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A17_ctrl_translator:uav_address
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A17_ctrl_translator:uav_write
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A17_ctrl_translator:uav_lock
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A17_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A17_ctrl_translator:uav_readdata -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A17_ctrl_translator:uav_readdatavalid -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A17_ctrl_translator:uav_debugaccess
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A17_ctrl_translator:uav_byteenable
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_B8_ctrl_translator:uav_waitrequest -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B8_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B8_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B8_ctrl_translator:uav_address
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B8_ctrl_translator:uav_write
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B8_ctrl_translator:uav_lock
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B8_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_B8_ctrl_translator:uav_readdata -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_B8_ctrl_translator:uav_readdatavalid -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B8_ctrl_translator:uav_debugaccess
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B8_ctrl_translator:uav_byteenable
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B24_ctrl_translator:uav_waitrequest -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B24_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B24_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B24_ctrl_translator:uav_address
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B24_ctrl_translator:uav_write
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B24_ctrl_translator:uav_lock
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B24_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B24_ctrl_translator:uav_readdata -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B24_ctrl_translator:uav_readdatavalid -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B24_ctrl_translator:uav_debugaccess
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B24_ctrl_translator:uav_byteenable
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_B7_ctrl_translator:uav_waitrequest -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B7_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B7_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B7_ctrl_translator:uav_address
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B7_ctrl_translator:uav_write
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B7_ctrl_translator:uav_lock
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B7_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_B7_ctrl_translator:uav_readdata -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_B7_ctrl_translator:uav_readdatavalid -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B7_ctrl_translator:uav_debugaccess
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B7_ctrl_translator:uav_byteenable
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B20_ctrl_translator:uav_waitrequest -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B20_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B20_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B20_ctrl_translator:uav_address
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B20_ctrl_translator:uav_write
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B20_ctrl_translator:uav_lock
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B20_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B20_ctrl_translator:uav_readdata -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B20_ctrl_translator:uav_readdatavalid -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B20_ctrl_translator:uav_debugaccess
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B20_ctrl_translator:uav_byteenable
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sam9_m1_translator_avalon_universal_master_0_waitrequest;                                // SAM9_M1_translator_avalon_universal_master_0_agent:av_waitrequest -> SAM9_M1_translator:uav_waitrequest
	wire   [2:0] sam9_m1_translator_avalon_universal_master_0_burstcount;                                 // SAM9_M1_translator:uav_burstcount -> SAM9_M1_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] sam9_m1_translator_avalon_universal_master_0_writedata;                                  // SAM9_M1_translator:uav_writedata -> SAM9_M1_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] sam9_m1_translator_avalon_universal_master_0_address;                                    // SAM9_M1_translator:uav_address -> SAM9_M1_translator_avalon_universal_master_0_agent:av_address
	wire         sam9_m1_translator_avalon_universal_master_0_lock;                                       // SAM9_M1_translator:uav_lock -> SAM9_M1_translator_avalon_universal_master_0_agent:av_lock
	wire         sam9_m1_translator_avalon_universal_master_0_write;                                      // SAM9_M1_translator:uav_write -> SAM9_M1_translator_avalon_universal_master_0_agent:av_write
	wire         sam9_m1_translator_avalon_universal_master_0_read;                                       // SAM9_M1_translator:uav_read -> SAM9_M1_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] sam9_m1_translator_avalon_universal_master_0_readdata;                                   // SAM9_M1_translator_avalon_universal_master_0_agent:av_readdata -> SAM9_M1_translator:uav_readdata
	wire         sam9_m1_translator_avalon_universal_master_0_debugaccess;                                // SAM9_M1_translator:uav_debugaccess -> SAM9_M1_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] sam9_m1_translator_avalon_universal_master_0_byteenable;                                 // SAM9_M1_translator:uav_byteenable -> SAM9_M1_translator_avalon_universal_master_0_agent:av_byteenable
	wire         sam9_m1_translator_avalon_universal_master_0_readdatavalid;                              // SAM9_M1_translator_avalon_universal_master_0_agent:av_readdatavalid -> SAM9_M1_translator:uav_readdatavalid
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A24_ctrl_translator:uav_waitrequest -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A24_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A24_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A24_ctrl_translator:uav_address
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A24_ctrl_translator:uav_write
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A24_ctrl_translator:uav_lock
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A24_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A24_ctrl_translator:uav_readdata -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A24_ctrl_translator:uav_readdatavalid -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A24_ctrl_translator:uav_debugaccess
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A24_ctrl_translator:uav_byteenable
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B16_ctrl_translator:uav_waitrequest -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B16_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B16_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B16_ctrl_translator:uav_address
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B16_ctrl_translator:uav_write
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B16_ctrl_translator:uav_lock
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B16_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B16_ctrl_translator:uav_readdata -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B16_ctrl_translator:uav_readdatavalid -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B16_ctrl_translator:uav_debugaccess
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B16_ctrl_translator:uav_byteenable
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A25_ctrl_translator:uav_waitrequest -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A25_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A25_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A25_ctrl_translator:uav_address
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A25_ctrl_translator:uav_write
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A25_ctrl_translator:uav_lock
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A25_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A25_ctrl_translator:uav_readdata -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A25_ctrl_translator:uav_readdatavalid -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A25_ctrl_translator:uav_debugaccess
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A25_ctrl_translator:uav_byteenable
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B15_ctrl_translator:uav_waitrequest -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B15_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B15_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B15_ctrl_translator:uav_address
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B15_ctrl_translator:uav_write
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B15_ctrl_translator:uav_lock
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B15_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B15_ctrl_translator:uav_readdata -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B15_ctrl_translator:uav_readdatavalid -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B15_ctrl_translator:uav_debugaccess
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B15_ctrl_translator:uav_byteenable
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_A7_ctrl_translator:uav_waitrequest -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A7_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A7_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A7_ctrl_translator:uav_address
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A7_ctrl_translator:uav_write
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A7_ctrl_translator:uav_lock
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A7_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_A7_ctrl_translator:uav_readdata -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_A7_ctrl_translator:uav_readdatavalid -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A7_ctrl_translator:uav_debugaccess
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A7_ctrl_translator:uav_byteenable
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B21_ctrl_translator:uav_waitrequest -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B21_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B21_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B21_ctrl_translator:uav_address
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B21_ctrl_translator:uav_write
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B21_ctrl_translator:uav_lock
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B21_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B21_ctrl_translator:uav_readdata -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B21_ctrl_translator:uav_readdatavalid -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B21_ctrl_translator:uav_debugaccess
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B21_ctrl_translator:uav_byteenable
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_A3_ctrl_translator:uav_waitrequest -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A3_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A3_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A3_ctrl_translator:uav_address
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A3_ctrl_translator:uav_write
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A3_ctrl_translator:uav_lock
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A3_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_A3_ctrl_translator:uav_readdata -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_A3_ctrl_translator:uav_readdatavalid -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A3_ctrl_translator:uav_debugaccess
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A3_ctrl_translator:uav_byteenable
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_B5_ctrl_translator:uav_waitrequest -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B5_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B5_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B5_ctrl_translator:uav_address
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B5_ctrl_translator:uav_write
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B5_ctrl_translator:uav_lock
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B5_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_B5_ctrl_translator:uav_readdata -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_B5_ctrl_translator:uav_readdatavalid -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B5_ctrl_translator:uav_debugaccess
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B5_ctrl_translator:uav_byteenable
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A14_ctrl_translator:uav_waitrequest -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A14_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A14_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A14_ctrl_translator:uav_address
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A14_ctrl_translator:uav_write
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A14_ctrl_translator:uav_lock
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A14_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A14_ctrl_translator:uav_readdata -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A14_ctrl_translator:uav_readdatavalid -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A14_ctrl_translator:uav_debugaccess
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A14_ctrl_translator:uav_byteenable
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B10_ctrl_translator:uav_waitrequest -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B10_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B10_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B10_ctrl_translator:uav_address
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B10_ctrl_translator:uav_write
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B10_ctrl_translator:uav_lock
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B10_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B10_ctrl_translator:uav_readdata -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B10_ctrl_translator:uav_readdatavalid -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B10_ctrl_translator:uav_debugaccess
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B10_ctrl_translator:uav_byteenable
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // FuncLED_1_LEDD_translator:uav_waitrequest -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> FuncLED_1_LEDD_translator:uav_burstcount
	wire  [31:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                   // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> FuncLED_1_LEDD_translator:uav_writedata
	wire  [31:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_address;                     // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> FuncLED_1_LEDD_translator:uav_address
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_write;                       // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> FuncLED_1_LEDD_translator:uav_write
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                        // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> FuncLED_1_LEDD_translator:uav_lock
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_read;                        // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> FuncLED_1_LEDD_translator:uav_read
	wire  [31:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                    // FuncLED_1_LEDD_translator:uav_readdata -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // FuncLED_1_LEDD_translator:uav_readdatavalid -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FuncLED_1_LEDD_translator:uav_debugaccess
	wire   [3:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> FuncLED_1_LEDD_translator:uav_byteenable
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;                // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                 // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;                // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B12_ctrl_translator:uav_waitrequest -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B12_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B12_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B12_ctrl_translator:uav_address
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B12_ctrl_translator:uav_write
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B12_ctrl_translator:uav_lock
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B12_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B12_ctrl_translator:uav_readdata -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B12_ctrl_translator:uav_readdatavalid -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B12_ctrl_translator:uav_debugaccess
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B12_ctrl_translator:uav_byteenable
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B14_ctrl_translator:uav_waitrequest -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B14_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B14_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B14_ctrl_translator:uav_address
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B14_ctrl_translator:uav_write
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B14_ctrl_translator:uav_lock
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B14_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B14_ctrl_translator:uav_readdata -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B14_ctrl_translator:uav_readdatavalid -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B14_ctrl_translator:uav_debugaccess
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B14_ctrl_translator:uav_byteenable
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_B6_ctrl_translator:uav_waitrequest -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B6_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B6_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B6_ctrl_translator:uav_address
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B6_ctrl_translator:uav_write
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B6_ctrl_translator:uav_lock
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B6_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_B6_ctrl_translator:uav_readdata -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_B6_ctrl_translator:uav_readdatavalid -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B6_ctrl_translator:uav_debugaccess
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B6_ctrl_translator:uav_byteenable
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_B9_ctrl_translator:uav_waitrequest -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B9_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B9_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B9_ctrl_translator:uav_address
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B9_ctrl_translator:uav_write
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B9_ctrl_translator:uav_lock
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B9_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_B9_ctrl_translator:uav_readdata -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_B9_ctrl_translator:uav_readdatavalid -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B9_ctrl_translator:uav_debugaccess
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B9_ctrl_translator:uav_byteenable
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A22_ctrl_translator:uav_waitrequest -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A22_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A22_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A22_ctrl_translator:uav_address
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A22_ctrl_translator:uav_write
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A22_ctrl_translator:uav_lock
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A22_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A22_ctrl_translator:uav_readdata -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A22_ctrl_translator:uav_readdatavalid -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A22_ctrl_translator:uav_debugaccess
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A22_ctrl_translator:uav_byteenable
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B23_ctrl_translator:uav_waitrequest -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B23_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B23_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B23_ctrl_translator:uav_address
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B23_ctrl_translator:uav_write
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B23_ctrl_translator:uav_lock
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B23_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B23_ctrl_translator:uav_readdata -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B23_ctrl_translator:uav_readdatavalid -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B23_ctrl_translator:uav_debugaccess
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B23_ctrl_translator:uav_byteenable
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B13_ctrl_translator:uav_waitrequest -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B13_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B13_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B13_ctrl_translator:uav_address
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B13_ctrl_translator:uav_write
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B13_ctrl_translator:uav_lock
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B13_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B13_ctrl_translator:uav_readdata -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B13_ctrl_translator:uav_readdatavalid -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B13_ctrl_translator:uav_debugaccess
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B13_ctrl_translator:uav_byteenable
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B25_ctrl_translator:uav_waitrequest -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B25_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B25_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B25_ctrl_translator:uav_address
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B25_ctrl_translator:uav_write
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B25_ctrl_translator:uav_lock
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B25_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B25_ctrl_translator:uav_readdata -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B25_ctrl_translator:uav_readdatavalid -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B25_ctrl_translator:uav_debugaccess
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B25_ctrl_translator:uav_byteenable
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A21_ctrl_translator:uav_waitrequest -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A21_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A21_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A21_ctrl_translator:uav_address
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A21_ctrl_translator:uav_write
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A21_ctrl_translator:uav_lock
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A21_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A21_ctrl_translator:uav_readdata -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A21_ctrl_translator:uav_readdatavalid -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A21_ctrl_translator:uav_debugaccess
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A21_ctrl_translator:uav_byteenable
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B18_ctrl_translator:uav_waitrequest -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B18_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B18_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B18_ctrl_translator:uav_address
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B18_ctrl_translator:uav_write
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B18_ctrl_translator:uav_lock
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B18_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B18_ctrl_translator:uav_readdata -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B18_ctrl_translator:uav_readdatavalid -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B18_ctrl_translator:uav_debugaccess
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B18_ctrl_translator:uav_byteenable
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shield_Admin_Ctrl_translator:uav_waitrequest -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shield_Admin_Ctrl_translator:uav_burstcount
	wire  [31:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shield_Admin_Ctrl_translator:uav_writedata
	wire  [31:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shield_Admin_Ctrl_translator:uav_address
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shield_Admin_Ctrl_translator:uav_write
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shield_Admin_Ctrl_translator:uav_lock
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shield_Admin_Ctrl_translator:uav_read
	wire  [31:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shield_Admin_Ctrl_translator:uav_readdata -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shield_Admin_Ctrl_translator:uav_readdatavalid -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shield_Admin_Ctrl_translator:uav_debugaccess
	wire   [3:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shield_Admin_Ctrl_translator:uav_byteenable
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B22_ctrl_translator:uav_waitrequest -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B22_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B22_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B22_ctrl_translator:uav_address
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B22_ctrl_translator:uav_write
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B22_ctrl_translator:uav_lock
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B22_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B22_ctrl_translator:uav_readdata -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B22_ctrl_translator:uav_readdatavalid -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B22_ctrl_translator:uav_debugaccess
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B22_ctrl_translator:uav_byteenable
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // SysID_SysID_translator:uav_waitrequest -> SysID_SysID_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_burstcount -> SysID_SysID_translator:uav_burstcount
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_writedata;                      // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_writedata -> SysID_SysID_translator:uav_writedata
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_address;                        // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_address -> SysID_SysID_translator:uav_address
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_write;                          // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_write -> SysID_SysID_translator:uav_write
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_lock;                           // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_lock -> SysID_SysID_translator:uav_lock
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_read;                           // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_read -> SysID_SysID_translator:uav_read
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdata;                       // SysID_SysID_translator:uav_readdata -> SysID_SysID_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // SysID_SysID_translator:uav_readdatavalid -> SysID_SysID_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SysID_SysID_translator:uav_debugaccess
	wire   [3:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_byteenable -> SysID_SysID_translator:uav_byteenable
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_data;                    // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_data -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A15_ctrl_translator:uav_waitrequest -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A15_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A15_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A15_ctrl_translator:uav_address
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A15_ctrl_translator:uav_write
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A15_ctrl_translator:uav_lock
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A15_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A15_ctrl_translator:uav_readdata -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A15_ctrl_translator:uav_readdatavalid -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A15_ctrl_translator:uav_debugaccess
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A15_ctrl_translator:uav_byteenable
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_B4_ctrl_translator:uav_waitrequest -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B4_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B4_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B4_ctrl_translator:uav_address
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B4_ctrl_translator:uav_write
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B4_ctrl_translator:uav_lock
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B4_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_B4_ctrl_translator:uav_readdata -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_B4_ctrl_translator:uav_readdatavalid -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B4_ctrl_translator:uav_debugaccess
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B4_ctrl_translator:uav_byteenable
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_A9_ctrl_translator:uav_waitrequest -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A9_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A9_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A9_ctrl_translator:uav_address
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A9_ctrl_translator:uav_write
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A9_ctrl_translator:uav_lock
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A9_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_A9_ctrl_translator:uav_readdata -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_A9_ctrl_translator:uav_readdatavalid -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A9_ctrl_translator:uav_debugaccess
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A9_ctrl_translator:uav_byteenable
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // FuncLED_3_LEDD_translator:uav_waitrequest -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> FuncLED_3_LEDD_translator:uav_burstcount
	wire  [31:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                   // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> FuncLED_3_LEDD_translator:uav_writedata
	wire  [31:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_address;                     // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> FuncLED_3_LEDD_translator:uav_address
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_write;                       // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> FuncLED_3_LEDD_translator:uav_write
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                        // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> FuncLED_3_LEDD_translator:uav_lock
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_read;                        // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> FuncLED_3_LEDD_translator:uav_read
	wire  [31:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                    // FuncLED_3_LEDD_translator:uav_readdata -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // FuncLED_3_LEDD_translator:uav_readdatavalid -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FuncLED_3_LEDD_translator:uav_debugaccess
	wire   [3:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> FuncLED_3_LEDD_translator:uav_byteenable
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;                // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                 // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;                // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_A8_ctrl_translator:uav_waitrequest -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A8_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A8_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A8_ctrl_translator:uav_address
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A8_ctrl_translator:uav_write
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A8_ctrl_translator:uav_lock
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A8_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_A8_ctrl_translator:uav_readdata -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_A8_ctrl_translator:uav_readdatavalid -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A8_ctrl_translator:uav_debugaccess
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A8_ctrl_translator:uav_byteenable
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_B3_ctrl_translator:uav_waitrequest -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B3_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B3_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B3_ctrl_translator:uav_address
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B3_ctrl_translator:uav_write
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B3_ctrl_translator:uav_lock
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B3_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_B3_ctrl_translator:uav_readdata -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_B3_ctrl_translator:uav_readdatavalid -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B3_ctrl_translator:uav_debugaccess
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B3_ctrl_translator:uav_byteenable
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_B17_ctrl_translator:uav_waitrequest -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_B17_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_B17_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_B17_ctrl_translator:uav_address
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_B17_ctrl_translator:uav_write
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_B17_ctrl_translator:uav_lock
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_B17_ctrl_translator:uav_read
	wire   [7:0] shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_B17_ctrl_translator:uav_readdata -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_B17_ctrl_translator:uav_readdatavalid -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_B17_ctrl_translator:uav_debugaccess
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_B17_ctrl_translator:uav_byteenable
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A13_ctrl_translator:uav_waitrequest -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A13_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A13_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A13_ctrl_translator:uav_address
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A13_ctrl_translator:uav_write
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A13_ctrl_translator:uav_lock
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A13_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A13_ctrl_translator:uav_readdata -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A13_ctrl_translator:uav_readdatavalid -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A13_ctrl_translator:uav_debugaccess
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A13_ctrl_translator:uav_byteenable
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A16_ctrl_translator:uav_waitrequest -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A16_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A16_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A16_ctrl_translator:uav_address
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A16_ctrl_translator:uav_write
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A16_ctrl_translator:uav_lock
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A16_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A16_ctrl_translator:uav_readdata -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A16_ctrl_translator:uav_readdatavalid -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A16_ctrl_translator:uav_debugaccess
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A16_ctrl_translator:uav_byteenable
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_A2_ctrl_translator:uav_waitrequest -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A2_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A2_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A2_ctrl_translator:uav_address
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A2_ctrl_translator:uav_write
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A2_ctrl_translator:uav_lock
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A2_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_A2_ctrl_translator:uav_readdata -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_A2_ctrl_translator:uav_readdatavalid -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A2_ctrl_translator:uav_debugaccess
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A2_ctrl_translator:uav_byteenable
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // FuncLED_2_LEDD_translator:uav_waitrequest -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> FuncLED_2_LEDD_translator:uav_burstcount
	wire  [31:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                   // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> FuncLED_2_LEDD_translator:uav_writedata
	wire  [31:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_address;                     // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> FuncLED_2_LEDD_translator:uav_address
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_write;                       // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> FuncLED_2_LEDD_translator:uav_write
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                        // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> FuncLED_2_LEDD_translator:uav_lock
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_read;                        // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> FuncLED_2_LEDD_translator:uav_read
	wire  [31:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                    // FuncLED_2_LEDD_translator:uav_readdata -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // FuncLED_2_LEDD_translator:uav_readdatavalid -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FuncLED_2_LEDD_translator:uav_debugaccess
	wire   [3:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> FuncLED_2_LEDD_translator:uav_byteenable
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;                // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                 // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;                // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // Shiled_IO_A5_ctrl_translator:uav_waitrequest -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A5_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;                // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A5_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                  // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A5_ctrl_translator:uav_address
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                    // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A5_ctrl_translator:uav_write
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                     // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A5_ctrl_translator:uav_lock
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                     // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A5_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // Shiled_IO_A5_ctrl_translator:uav_readdata -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // Shiled_IO_A5_ctrl_translator:uav_readdatavalid -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A5_ctrl_translator:uav_debugaccess
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A5_ctrl_translator:uav_byteenable
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;              // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A23_ctrl_translator:uav_waitrequest -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A23_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A23_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A23_ctrl_translator:uav_address
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A23_ctrl_translator:uav_write
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A23_ctrl_translator:uav_lock
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A23_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A23_ctrl_translator:uav_readdata -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A23_ctrl_translator:uav_readdatavalid -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A23_ctrl_translator:uav_debugaccess
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A23_ctrl_translator:uav_byteenable
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shiled_IO_A18_ctrl_translator:uav_waitrequest -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shiled_IO_A18_ctrl_translator:uav_burstcount
	wire   [7:0] shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shiled_IO_A18_ctrl_translator:uav_writedata
	wire  [31:0] shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shiled_IO_A18_ctrl_translator:uav_address
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shiled_IO_A18_ctrl_translator:uav_write
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shiled_IO_A18_ctrl_translator:uav_lock
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shiled_IO_A18_ctrl_translator:uav_read
	wire   [7:0] shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shiled_IO_A18_ctrl_translator:uav_readdata -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shiled_IO_A18_ctrl_translator:uav_readdatavalid -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shiled_IO_A18_ctrl_translator:uav_debugaccess
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shiled_IO_A18_ctrl_translator:uav_byteenable
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [66:0] shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [66:0] shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [7:0] shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sam9_m1_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // SAM9_M1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         sam9_m1_translator_avalon_universal_master_0_agent_cp_valid;                             // SAM9_M1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         sam9_m1_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // SAM9_M1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [92:0] sam9_m1_translator_avalon_universal_master_0_agent_cp_data;                              // SAM9_M1_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         sam9_m1_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router:sink_ready -> SAM9_M1_translator_avalon_universal_master_0_agent:cp_ready
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_valid;                          // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [92:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rp_data;                           // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router:sink_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent:rp_ready
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                       // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [92:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_data;                        // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_001:sink_ready -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                       // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [92:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_data;                        // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_002:sink_ready -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                       // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [92:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_data;                        // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_003:sink_ready -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                       // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [92:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_data;                        // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_004:sink_ready -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [92:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_005:sink_ready -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [65:0] shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_006:sink_ready -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [65:0] shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_007:sink_ready -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [65:0] shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_008:sink_ready -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [65:0] shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_009:sink_ready -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [65:0] shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_010:sink_ready -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [65:0] shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_011:sink_ready -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [65:0] shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_012:sink_ready -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [65:0] shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_013:sink_ready -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [65:0] shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire         shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_014:sink_ready -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [65:0] shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire         shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_015:sink_ready -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [65:0] shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire         shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_016:sink_ready -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [65:0] shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire         shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_017:sink_ready -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [65:0] shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire         shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_018:sink_ready -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [65:0] shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire         shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_019:sink_ready -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [65:0] shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire         shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_020:sink_ready -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [65:0] shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire         shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_021:sink_ready -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire  [65:0] shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire         shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_022:sink_ready -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire  [65:0] shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire         shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_023:sink_ready -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire  [65:0] shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire         shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_024:sink_ready -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire  [65:0] shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire         shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_025:sink_ready -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	wire  [65:0] shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	wire         shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_026:sink_ready -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	wire  [65:0] shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	wire         shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_027:sink_ready -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	wire  [65:0] shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	wire         shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_028:sink_ready -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_029:sink_endofpacket
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_029:sink_valid
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_029:sink_startofpacket
	wire  [65:0] shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_029:sink_data
	wire         shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_029:sink_ready -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_030:sink_endofpacket
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_030:sink_valid
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_030:sink_startofpacket
	wire  [65:0] shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_030:sink_data
	wire         shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_030:sink_ready -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_031:sink_endofpacket
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_031:sink_valid
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_031:sink_startofpacket
	wire  [65:0] shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_031:sink_data
	wire         shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_031:sink_ready -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_032:sink_endofpacket
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_032:sink_valid
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_032:sink_startofpacket
	wire  [65:0] shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_032:sink_data
	wire         shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_032:sink_ready -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_033:sink_endofpacket
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_033:sink_valid
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_033:sink_startofpacket
	wire  [65:0] shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_033:sink_data
	wire         shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_033:sink_ready -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_034:sink_endofpacket
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_034:sink_valid
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_034:sink_startofpacket
	wire  [65:0] shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_034:sink_data
	wire         shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_034:sink_ready -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_035:sink_endofpacket
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_035:sink_valid
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_035:sink_startofpacket
	wire  [65:0] shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_035:sink_data
	wire         shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_035:sink_ready -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_036:sink_endofpacket
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_036:sink_valid
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_036:sink_startofpacket
	wire  [65:0] shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_036:sink_data
	wire         shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_036:sink_ready -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_037:sink_endofpacket
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_037:sink_valid
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_037:sink_startofpacket
	wire  [65:0] shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_037:sink_data
	wire         shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_037:sink_ready -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_038:sink_endofpacket
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_038:sink_valid
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_038:sink_startofpacket
	wire  [65:0] shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_038:sink_data
	wire         shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_038:sink_ready -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_039:sink_endofpacket
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_039:sink_valid
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_039:sink_startofpacket
	wire  [65:0] shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_039:sink_data
	wire         shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_039:sink_ready -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_040:sink_endofpacket
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_040:sink_valid
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_040:sink_startofpacket
	wire  [65:0] shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_040:sink_data
	wire         shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_040:sink_ready -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_041:sink_endofpacket
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                    // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_041:sink_valid
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_041:sink_startofpacket
	wire  [65:0] shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                     // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_041:sink_data
	wire         shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_041:sink_ready -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_042:sink_endofpacket
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_042:sink_valid
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_042:sink_startofpacket
	wire  [65:0] shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_042:sink_data
	wire         shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_042:sink_ready -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_043:sink_endofpacket
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_043:sink_valid
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_043:sink_startofpacket
	wire  [65:0] shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_043:sink_data
	wire         shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_043:sink_ready -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_044:sink_endofpacket
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_044:sink_valid
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_044:sink_startofpacket
	wire  [65:0] shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_044:sink_data
	wire         shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_044:sink_ready -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_045:sink_endofpacket
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_045:sink_valid
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_045:sink_startofpacket
	wire  [65:0] shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_045:sink_data
	wire         shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_045:sink_ready -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_046:sink_endofpacket
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_046:sink_valid
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_046:sink_startofpacket
	wire  [65:0] shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_046:sink_data
	wire         shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_046:sink_ready -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_047:sink_endofpacket
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_047:sink_valid
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_047:sink_startofpacket
	wire  [65:0] shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_047:sink_data
	wire         shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_047:sink_ready -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_048:sink_endofpacket
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_048:sink_valid
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_048:sink_startofpacket
	wire  [65:0] shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_048:sink_data
	wire         shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_048:sink_ready -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_049:sink_endofpacket
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_049:sink_valid
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_049:sink_startofpacket
	wire  [65:0] shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_049:sink_data
	wire         shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_049:sink_ready -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_050:sink_endofpacket
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_050:sink_valid
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_050:sink_startofpacket
	wire  [65:0] shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_050:sink_data
	wire         shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_050:sink_ready -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_051:sink_endofpacket
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_051:sink_valid
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_051:sink_startofpacket
	wire  [65:0] shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_051:sink_data
	wire         shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_051:sink_ready -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_052:sink_endofpacket
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_052:sink_valid
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_052:sink_startofpacket
	wire  [65:0] shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_052:sink_data
	wire         shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_052:sink_ready -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_053:sink_endofpacket
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_053:sink_valid
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_053:sink_startofpacket
	wire  [65:0] shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_053:sink_data
	wire         shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_053:sink_ready -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_054:sink_endofpacket
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_054:sink_valid
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_054:sink_startofpacket
	wire  [65:0] shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_054:sink_data
	wire         shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_054:sink_ready -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_055:sink_endofpacket
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_055:sink_valid
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_055:sink_startofpacket
	wire  [65:0] shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_055:sink_data
	wire         shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_055:sink_ready -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_056:sink_endofpacket
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_056:sink_valid
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_056:sink_startofpacket
	wire  [65:0] shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_056:sink_data
	wire         shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_056:sink_ready -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_057:sink_endofpacket
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_057:sink_valid
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_057:sink_startofpacket
	wire  [65:0] shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_057:sink_data
	wire         shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_057:sink_ready -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                             // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                   // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                           // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [92:0] addr_router_src_data;                                                                    // addr_router:src_data -> limiter:cmd_sink_data
	wire  [57:0] addr_router_src_channel;                                                                 // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                   // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                             // limiter:rsp_src_endofpacket -> SAM9_M1_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                   // limiter:rsp_src_valid -> SAM9_M1_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                           // limiter:rsp_src_startofpacket -> SAM9_M1_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [92:0] limiter_rsp_src_data;                                                                    // limiter:rsp_src_data -> SAM9_M1_translator_avalon_universal_master_0_agent:rp_data
	wire  [57:0] limiter_rsp_src_channel;                                                                 // limiter:rsp_src_channel -> SAM9_M1_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                   // SAM9_M1_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         burst_adapter_source0_endofpacket;                                                       // burst_adapter:source0_endofpacket -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                             // burst_adapter:source0_valid -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                     // burst_adapter:source0_startofpacket -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_source0_data;                                                              // burst_adapter:source0_data -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                             // Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire  [57:0] burst_adapter_source0_channel;                                                           // burst_adapter:source0_channel -> Shiled_IO_B0_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_001_source0_endofpacket;                                                   // burst_adapter_001:source0_endofpacket -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_001_source0_valid;                                                         // burst_adapter_001:source0_valid -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_001_source0_startofpacket;                                                 // burst_adapter_001:source0_startofpacket -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_001_source0_data;                                                          // burst_adapter_001:source0_data -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_001_source0_ready;                                                         // Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire  [57:0] burst_adapter_001_source0_channel;                                                       // burst_adapter_001:source0_channel -> Shiled_IO_B2_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_002_source0_endofpacket;                                                   // burst_adapter_002:source0_endofpacket -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_002_source0_valid;                                                         // burst_adapter_002:source0_valid -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_002_source0_startofpacket;                                                 // burst_adapter_002:source0_startofpacket -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_002_source0_data;                                                          // burst_adapter_002:source0_data -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_002_source0_ready;                                                         // Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire  [57:0] burst_adapter_002_source0_channel;                                                       // burst_adapter_002:source0_channel -> Shiled_IO_A12_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_003_source0_endofpacket;                                                   // burst_adapter_003:source0_endofpacket -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_003_source0_valid;                                                         // burst_adapter_003:source0_valid -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_003_source0_startofpacket;                                                 // burst_adapter_003:source0_startofpacket -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_003_source0_data;                                                          // burst_adapter_003:source0_data -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_003_source0_ready;                                                         // Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire  [57:0] burst_adapter_003_source0_channel;                                                       // burst_adapter_003:source0_channel -> Shiled_IO_A11_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_004_source0_endofpacket;                                                   // burst_adapter_004:source0_endofpacket -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_004_source0_valid;                                                         // burst_adapter_004:source0_valid -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_004_source0_startofpacket;                                                 // burst_adapter_004:source0_startofpacket -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_004_source0_data;                                                          // burst_adapter_004:source0_data -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_004_source0_ready;                                                         // Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_004:source0_ready
	wire  [57:0] burst_adapter_004_source0_channel;                                                       // burst_adapter_004:source0_channel -> Shiled_IO_A1_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_005_source0_endofpacket;                                                   // burst_adapter_005:source0_endofpacket -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_005_source0_valid;                                                         // burst_adapter_005:source0_valid -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_005_source0_startofpacket;                                                 // burst_adapter_005:source0_startofpacket -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_005_source0_data;                                                          // burst_adapter_005:source0_data -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_005_source0_ready;                                                         // Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_005:source0_ready
	wire  [57:0] burst_adapter_005_source0_channel;                                                       // burst_adapter_005:source0_channel -> Shiled_IO_A0_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_006_source0_endofpacket;                                                   // burst_adapter_006:source0_endofpacket -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_006_source0_valid;                                                         // burst_adapter_006:source0_valid -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_006_source0_startofpacket;                                                 // burst_adapter_006:source0_startofpacket -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_006_source0_data;                                                          // burst_adapter_006:source0_data -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_006_source0_ready;                                                         // Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_006:source0_ready
	wire  [57:0] burst_adapter_006_source0_channel;                                                       // burst_adapter_006:source0_channel -> Shiled_IO_B19_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_007_source0_endofpacket;                                                   // burst_adapter_007:source0_endofpacket -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_007_source0_valid;                                                         // burst_adapter_007:source0_valid -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_007_source0_startofpacket;                                                 // burst_adapter_007:source0_startofpacket -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_007_source0_data;                                                          // burst_adapter_007:source0_data -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_007_source0_ready;                                                         // Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_007:source0_ready
	wire  [57:0] burst_adapter_007_source0_channel;                                                       // burst_adapter_007:source0_channel -> Shiled_IO_A10_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_008_source0_endofpacket;                                                   // burst_adapter_008:source0_endofpacket -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_008_source0_valid;                                                         // burst_adapter_008:source0_valid -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_008_source0_startofpacket;                                                 // burst_adapter_008:source0_startofpacket -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_008_source0_data;                                                          // burst_adapter_008:source0_data -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_008_source0_ready;                                                         // Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_008:source0_ready
	wire  [57:0] burst_adapter_008_source0_channel;                                                       // burst_adapter_008:source0_channel -> Shiled_IO_A19_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_009_source0_endofpacket;                                                   // burst_adapter_009:source0_endofpacket -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_009_source0_valid;                                                         // burst_adapter_009:source0_valid -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_009_source0_startofpacket;                                                 // burst_adapter_009:source0_startofpacket -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_009_source0_data;                                                          // burst_adapter_009:source0_data -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_009_source0_ready;                                                         // Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_009:source0_ready
	wire  [57:0] burst_adapter_009_source0_channel;                                                       // burst_adapter_009:source0_channel -> Shiled_IO_B1_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_010_source0_endofpacket;                                                   // burst_adapter_010:source0_endofpacket -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_010_source0_valid;                                                         // burst_adapter_010:source0_valid -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_010_source0_startofpacket;                                                 // burst_adapter_010:source0_startofpacket -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_010_source0_data;                                                          // burst_adapter_010:source0_data -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_010_source0_ready;                                                         // Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_010:source0_ready
	wire  [57:0] burst_adapter_010_source0_channel;                                                       // burst_adapter_010:source0_channel -> Shiled_IO_A6_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_011_source0_endofpacket;                                                   // burst_adapter_011:source0_endofpacket -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_011_source0_valid;                                                         // burst_adapter_011:source0_valid -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_011_source0_startofpacket;                                                 // burst_adapter_011:source0_startofpacket -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_011_source0_data;                                                          // burst_adapter_011:source0_data -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_011_source0_ready;                                                         // Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_011:source0_ready
	wire  [57:0] burst_adapter_011_source0_channel;                                                       // burst_adapter_011:source0_channel -> Shiled_IO_A4_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_012_source0_endofpacket;                                                   // burst_adapter_012:source0_endofpacket -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_012_source0_valid;                                                         // burst_adapter_012:source0_valid -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_012_source0_startofpacket;                                                 // burst_adapter_012:source0_startofpacket -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_012_source0_data;                                                          // burst_adapter_012:source0_data -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_012_source0_ready;                                                         // Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_012:source0_ready
	wire  [57:0] burst_adapter_012_source0_channel;                                                       // burst_adapter_012:source0_channel -> Shiled_IO_A20_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_013_source0_endofpacket;                                                   // burst_adapter_013:source0_endofpacket -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_013_source0_valid;                                                         // burst_adapter_013:source0_valid -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_013_source0_startofpacket;                                                 // burst_adapter_013:source0_startofpacket -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_013_source0_data;                                                          // burst_adapter_013:source0_data -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_013_source0_ready;                                                         // Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_013:source0_ready
	wire  [57:0] burst_adapter_013_source0_channel;                                                       // burst_adapter_013:source0_channel -> Shiled_IO_B11_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_014_source0_endofpacket;                                                   // burst_adapter_014:source0_endofpacket -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_014_source0_valid;                                                         // burst_adapter_014:source0_valid -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_014_source0_startofpacket;                                                 // burst_adapter_014:source0_startofpacket -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_014_source0_data;                                                          // burst_adapter_014:source0_data -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_014_source0_ready;                                                         // Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_014:source0_ready
	wire  [57:0] burst_adapter_014_source0_channel;                                                       // burst_adapter_014:source0_channel -> Shiled_IO_A17_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_015_source0_endofpacket;                                                   // burst_adapter_015:source0_endofpacket -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_015_source0_valid;                                                         // burst_adapter_015:source0_valid -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_015_source0_startofpacket;                                                 // burst_adapter_015:source0_startofpacket -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_015_source0_data;                                                          // burst_adapter_015:source0_data -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_015_source0_ready;                                                         // Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_015:source0_ready
	wire  [57:0] burst_adapter_015_source0_channel;                                                       // burst_adapter_015:source0_channel -> Shiled_IO_B8_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_016_source0_endofpacket;                                                   // burst_adapter_016:source0_endofpacket -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_016_source0_valid;                                                         // burst_adapter_016:source0_valid -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_016_source0_startofpacket;                                                 // burst_adapter_016:source0_startofpacket -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_016_source0_data;                                                          // burst_adapter_016:source0_data -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_016_source0_ready;                                                         // Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_016:source0_ready
	wire  [57:0] burst_adapter_016_source0_channel;                                                       // burst_adapter_016:source0_channel -> Shiled_IO_B24_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_017_source0_endofpacket;                                                   // burst_adapter_017:source0_endofpacket -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_017_source0_valid;                                                         // burst_adapter_017:source0_valid -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_017_source0_startofpacket;                                                 // burst_adapter_017:source0_startofpacket -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_017_source0_data;                                                          // burst_adapter_017:source0_data -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_017_source0_ready;                                                         // Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_017:source0_ready
	wire  [57:0] burst_adapter_017_source0_channel;                                                       // burst_adapter_017:source0_channel -> Shiled_IO_B7_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_018_source0_endofpacket;                                                   // burst_adapter_018:source0_endofpacket -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_018_source0_valid;                                                         // burst_adapter_018:source0_valid -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_018_source0_startofpacket;                                                 // burst_adapter_018:source0_startofpacket -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_018_source0_data;                                                          // burst_adapter_018:source0_data -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_018_source0_ready;                                                         // Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_018:source0_ready
	wire  [57:0] burst_adapter_018_source0_channel;                                                       // burst_adapter_018:source0_channel -> Shiled_IO_B20_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_019_source0_endofpacket;                                                   // burst_adapter_019:source0_endofpacket -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_019_source0_valid;                                                         // burst_adapter_019:source0_valid -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_019_source0_startofpacket;                                                 // burst_adapter_019:source0_startofpacket -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_019_source0_data;                                                          // burst_adapter_019:source0_data -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_019_source0_ready;                                                         // Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_019:source0_ready
	wire  [57:0] burst_adapter_019_source0_channel;                                                       // burst_adapter_019:source0_channel -> Shiled_IO_A24_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_020_source0_endofpacket;                                                   // burst_adapter_020:source0_endofpacket -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_020_source0_valid;                                                         // burst_adapter_020:source0_valid -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_020_source0_startofpacket;                                                 // burst_adapter_020:source0_startofpacket -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_020_source0_data;                                                          // burst_adapter_020:source0_data -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_020_source0_ready;                                                         // Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_020:source0_ready
	wire  [57:0] burst_adapter_020_source0_channel;                                                       // burst_adapter_020:source0_channel -> Shiled_IO_B16_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_021_source0_endofpacket;                                                   // burst_adapter_021:source0_endofpacket -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_021_source0_valid;                                                         // burst_adapter_021:source0_valid -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_021_source0_startofpacket;                                                 // burst_adapter_021:source0_startofpacket -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_021_source0_data;                                                          // burst_adapter_021:source0_data -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_021_source0_ready;                                                         // Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_021:source0_ready
	wire  [57:0] burst_adapter_021_source0_channel;                                                       // burst_adapter_021:source0_channel -> Shiled_IO_A25_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_022_source0_endofpacket;                                                   // burst_adapter_022:source0_endofpacket -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_022_source0_valid;                                                         // burst_adapter_022:source0_valid -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_022_source0_startofpacket;                                                 // burst_adapter_022:source0_startofpacket -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_022_source0_data;                                                          // burst_adapter_022:source0_data -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_022_source0_ready;                                                         // Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_022:source0_ready
	wire  [57:0] burst_adapter_022_source0_channel;                                                       // burst_adapter_022:source0_channel -> Shiled_IO_B15_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_023_source0_endofpacket;                                                   // burst_adapter_023:source0_endofpacket -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_023_source0_valid;                                                         // burst_adapter_023:source0_valid -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_023_source0_startofpacket;                                                 // burst_adapter_023:source0_startofpacket -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_023_source0_data;                                                          // burst_adapter_023:source0_data -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_023_source0_ready;                                                         // Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_023:source0_ready
	wire  [57:0] burst_adapter_023_source0_channel;                                                       // burst_adapter_023:source0_channel -> Shiled_IO_A7_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_024_source0_endofpacket;                                                   // burst_adapter_024:source0_endofpacket -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_024_source0_valid;                                                         // burst_adapter_024:source0_valid -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_024_source0_startofpacket;                                                 // burst_adapter_024:source0_startofpacket -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_024_source0_data;                                                          // burst_adapter_024:source0_data -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_024_source0_ready;                                                         // Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_024:source0_ready
	wire  [57:0] burst_adapter_024_source0_channel;                                                       // burst_adapter_024:source0_channel -> Shiled_IO_B21_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_025_source0_endofpacket;                                                   // burst_adapter_025:source0_endofpacket -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_025_source0_valid;                                                         // burst_adapter_025:source0_valid -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_025_source0_startofpacket;                                                 // burst_adapter_025:source0_startofpacket -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_025_source0_data;                                                          // burst_adapter_025:source0_data -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_025_source0_ready;                                                         // Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_025:source0_ready
	wire  [57:0] burst_adapter_025_source0_channel;                                                       // burst_adapter_025:source0_channel -> Shiled_IO_A3_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_026_source0_endofpacket;                                                   // burst_adapter_026:source0_endofpacket -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_026_source0_valid;                                                         // burst_adapter_026:source0_valid -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_026_source0_startofpacket;                                                 // burst_adapter_026:source0_startofpacket -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_026_source0_data;                                                          // burst_adapter_026:source0_data -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_026_source0_ready;                                                         // Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_026:source0_ready
	wire  [57:0] burst_adapter_026_source0_channel;                                                       // burst_adapter_026:source0_channel -> Shiled_IO_B5_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_027_source0_endofpacket;                                                   // burst_adapter_027:source0_endofpacket -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_027_source0_valid;                                                         // burst_adapter_027:source0_valid -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_027_source0_startofpacket;                                                 // burst_adapter_027:source0_startofpacket -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_027_source0_data;                                                          // burst_adapter_027:source0_data -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_027_source0_ready;                                                         // Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_027:source0_ready
	wire  [57:0] burst_adapter_027_source0_channel;                                                       // burst_adapter_027:source0_channel -> Shiled_IO_A14_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_028_source0_endofpacket;                                                   // burst_adapter_028:source0_endofpacket -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_028_source0_valid;                                                         // burst_adapter_028:source0_valid -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_028_source0_startofpacket;                                                 // burst_adapter_028:source0_startofpacket -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_028_source0_data;                                                          // burst_adapter_028:source0_data -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_028_source0_ready;                                                         // Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_028:source0_ready
	wire  [57:0] burst_adapter_028_source0_channel;                                                       // burst_adapter_028:source0_channel -> Shiled_IO_B10_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_029_source0_endofpacket;                                                   // burst_adapter_029:source0_endofpacket -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_029_source0_valid;                                                         // burst_adapter_029:source0_valid -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_029_source0_startofpacket;                                                 // burst_adapter_029:source0_startofpacket -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_029_source0_data;                                                          // burst_adapter_029:source0_data -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_029_source0_ready;                                                         // Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_029:source0_ready
	wire  [57:0] burst_adapter_029_source0_channel;                                                       // burst_adapter_029:source0_channel -> Shiled_IO_B12_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_030_source0_endofpacket;                                                   // burst_adapter_030:source0_endofpacket -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_030_source0_valid;                                                         // burst_adapter_030:source0_valid -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_030_source0_startofpacket;                                                 // burst_adapter_030:source0_startofpacket -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_030_source0_data;                                                          // burst_adapter_030:source0_data -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_030_source0_ready;                                                         // Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_030:source0_ready
	wire  [57:0] burst_adapter_030_source0_channel;                                                       // burst_adapter_030:source0_channel -> Shiled_IO_B14_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_031_source0_endofpacket;                                                   // burst_adapter_031:source0_endofpacket -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_031_source0_valid;                                                         // burst_adapter_031:source0_valid -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_031_source0_startofpacket;                                                 // burst_adapter_031:source0_startofpacket -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_031_source0_data;                                                          // burst_adapter_031:source0_data -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_031_source0_ready;                                                         // Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_031:source0_ready
	wire  [57:0] burst_adapter_031_source0_channel;                                                       // burst_adapter_031:source0_channel -> Shiled_IO_B6_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_032_source0_endofpacket;                                                   // burst_adapter_032:source0_endofpacket -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_032_source0_valid;                                                         // burst_adapter_032:source0_valid -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_032_source0_startofpacket;                                                 // burst_adapter_032:source0_startofpacket -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_032_source0_data;                                                          // burst_adapter_032:source0_data -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_032_source0_ready;                                                         // Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_032:source0_ready
	wire  [57:0] burst_adapter_032_source0_channel;                                                       // burst_adapter_032:source0_channel -> Shiled_IO_B9_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_033_source0_endofpacket;                                                   // burst_adapter_033:source0_endofpacket -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_033_source0_valid;                                                         // burst_adapter_033:source0_valid -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_033_source0_startofpacket;                                                 // burst_adapter_033:source0_startofpacket -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_033_source0_data;                                                          // burst_adapter_033:source0_data -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_033_source0_ready;                                                         // Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_033:source0_ready
	wire  [57:0] burst_adapter_033_source0_channel;                                                       // burst_adapter_033:source0_channel -> Shiled_IO_A22_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_034_source0_endofpacket;                                                   // burst_adapter_034:source0_endofpacket -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_034_source0_valid;                                                         // burst_adapter_034:source0_valid -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_034_source0_startofpacket;                                                 // burst_adapter_034:source0_startofpacket -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_034_source0_data;                                                          // burst_adapter_034:source0_data -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_034_source0_ready;                                                         // Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_034:source0_ready
	wire  [57:0] burst_adapter_034_source0_channel;                                                       // burst_adapter_034:source0_channel -> Shiled_IO_B23_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_035_source0_endofpacket;                                                   // burst_adapter_035:source0_endofpacket -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_035_source0_valid;                                                         // burst_adapter_035:source0_valid -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_035_source0_startofpacket;                                                 // burst_adapter_035:source0_startofpacket -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_035_source0_data;                                                          // burst_adapter_035:source0_data -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_035_source0_ready;                                                         // Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_035:source0_ready
	wire  [57:0] burst_adapter_035_source0_channel;                                                       // burst_adapter_035:source0_channel -> Shiled_IO_B13_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_036_source0_endofpacket;                                                   // burst_adapter_036:source0_endofpacket -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_036_source0_valid;                                                         // burst_adapter_036:source0_valid -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_036_source0_startofpacket;                                                 // burst_adapter_036:source0_startofpacket -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_036_source0_data;                                                          // burst_adapter_036:source0_data -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_036_source0_ready;                                                         // Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_036:source0_ready
	wire  [57:0] burst_adapter_036_source0_channel;                                                       // burst_adapter_036:source0_channel -> Shiled_IO_B25_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_037_source0_endofpacket;                                                   // burst_adapter_037:source0_endofpacket -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_037_source0_valid;                                                         // burst_adapter_037:source0_valid -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_037_source0_startofpacket;                                                 // burst_adapter_037:source0_startofpacket -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_037_source0_data;                                                          // burst_adapter_037:source0_data -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_037_source0_ready;                                                         // Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_037:source0_ready
	wire  [57:0] burst_adapter_037_source0_channel;                                                       // burst_adapter_037:source0_channel -> Shiled_IO_A21_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_038_source0_endofpacket;                                                   // burst_adapter_038:source0_endofpacket -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_038_source0_valid;                                                         // burst_adapter_038:source0_valid -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_038_source0_startofpacket;                                                 // burst_adapter_038:source0_startofpacket -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_038_source0_data;                                                          // burst_adapter_038:source0_data -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_038_source0_ready;                                                         // Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_038:source0_ready
	wire  [57:0] burst_adapter_038_source0_channel;                                                       // burst_adapter_038:source0_channel -> Shiled_IO_B18_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_039_source0_endofpacket;                                                   // burst_adapter_039:source0_endofpacket -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_039_source0_valid;                                                         // burst_adapter_039:source0_valid -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_039_source0_startofpacket;                                                 // burst_adapter_039:source0_startofpacket -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_039_source0_data;                                                          // burst_adapter_039:source0_data -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_039_source0_ready;                                                         // Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_039:source0_ready
	wire  [57:0] burst_adapter_039_source0_channel;                                                       // burst_adapter_039:source0_channel -> Shiled_IO_B22_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_040_source0_endofpacket;                                                   // burst_adapter_040:source0_endofpacket -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_040_source0_valid;                                                         // burst_adapter_040:source0_valid -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_040_source0_startofpacket;                                                 // burst_adapter_040:source0_startofpacket -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_040_source0_data;                                                          // burst_adapter_040:source0_data -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_040_source0_ready;                                                         // Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_040:source0_ready
	wire  [57:0] burst_adapter_040_source0_channel;                                                       // burst_adapter_040:source0_channel -> Shiled_IO_A15_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_041_source0_endofpacket;                                                   // burst_adapter_041:source0_endofpacket -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_041_source0_valid;                                                         // burst_adapter_041:source0_valid -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_041_source0_startofpacket;                                                 // burst_adapter_041:source0_startofpacket -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_041_source0_data;                                                          // burst_adapter_041:source0_data -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_041_source0_ready;                                                         // Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_041:source0_ready
	wire  [57:0] burst_adapter_041_source0_channel;                                                       // burst_adapter_041:source0_channel -> Shiled_IO_B4_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_042_source0_endofpacket;                                                   // burst_adapter_042:source0_endofpacket -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_042_source0_valid;                                                         // burst_adapter_042:source0_valid -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_042_source0_startofpacket;                                                 // burst_adapter_042:source0_startofpacket -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_042_source0_data;                                                          // burst_adapter_042:source0_data -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_042_source0_ready;                                                         // Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_042:source0_ready
	wire  [57:0] burst_adapter_042_source0_channel;                                                       // burst_adapter_042:source0_channel -> Shiled_IO_A9_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_043_source0_endofpacket;                                                   // burst_adapter_043:source0_endofpacket -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_043_source0_valid;                                                         // burst_adapter_043:source0_valid -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_043_source0_startofpacket;                                                 // burst_adapter_043:source0_startofpacket -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_043_source0_data;                                                          // burst_adapter_043:source0_data -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_043_source0_ready;                                                         // Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_043:source0_ready
	wire  [57:0] burst_adapter_043_source0_channel;                                                       // burst_adapter_043:source0_channel -> Shiled_IO_A8_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_044_source0_endofpacket;                                                   // burst_adapter_044:source0_endofpacket -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_044_source0_valid;                                                         // burst_adapter_044:source0_valid -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_044_source0_startofpacket;                                                 // burst_adapter_044:source0_startofpacket -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_044_source0_data;                                                          // burst_adapter_044:source0_data -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_044_source0_ready;                                                         // Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_044:source0_ready
	wire  [57:0] burst_adapter_044_source0_channel;                                                       // burst_adapter_044:source0_channel -> Shiled_IO_B3_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_045_source0_endofpacket;                                                   // burst_adapter_045:source0_endofpacket -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_045_source0_valid;                                                         // burst_adapter_045:source0_valid -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_045_source0_startofpacket;                                                 // burst_adapter_045:source0_startofpacket -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_045_source0_data;                                                          // burst_adapter_045:source0_data -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_045_source0_ready;                                                         // Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_045:source0_ready
	wire  [57:0] burst_adapter_045_source0_channel;                                                       // burst_adapter_045:source0_channel -> Shiled_IO_B17_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_046_source0_endofpacket;                                                   // burst_adapter_046:source0_endofpacket -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_046_source0_valid;                                                         // burst_adapter_046:source0_valid -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_046_source0_startofpacket;                                                 // burst_adapter_046:source0_startofpacket -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_046_source0_data;                                                          // burst_adapter_046:source0_data -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_046_source0_ready;                                                         // Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_046:source0_ready
	wire  [57:0] burst_adapter_046_source0_channel;                                                       // burst_adapter_046:source0_channel -> Shiled_IO_A13_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_047_source0_endofpacket;                                                   // burst_adapter_047:source0_endofpacket -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_047_source0_valid;                                                         // burst_adapter_047:source0_valid -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_047_source0_startofpacket;                                                 // burst_adapter_047:source0_startofpacket -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_047_source0_data;                                                          // burst_adapter_047:source0_data -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_047_source0_ready;                                                         // Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_047:source0_ready
	wire  [57:0] burst_adapter_047_source0_channel;                                                       // burst_adapter_047:source0_channel -> Shiled_IO_A16_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_048_source0_endofpacket;                                                   // burst_adapter_048:source0_endofpacket -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_048_source0_valid;                                                         // burst_adapter_048:source0_valid -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_048_source0_startofpacket;                                                 // burst_adapter_048:source0_startofpacket -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_048_source0_data;                                                          // burst_adapter_048:source0_data -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_048_source0_ready;                                                         // Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_048:source0_ready
	wire  [57:0] burst_adapter_048_source0_channel;                                                       // burst_adapter_048:source0_channel -> Shiled_IO_A2_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_049_source0_endofpacket;                                                   // burst_adapter_049:source0_endofpacket -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_049_source0_valid;                                                         // burst_adapter_049:source0_valid -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_049_source0_startofpacket;                                                 // burst_adapter_049:source0_startofpacket -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_049_source0_data;                                                          // burst_adapter_049:source0_data -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_049_source0_ready;                                                         // Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_049:source0_ready
	wire  [57:0] burst_adapter_049_source0_channel;                                                       // burst_adapter_049:source0_channel -> Shiled_IO_A5_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_050_source0_endofpacket;                                                   // burst_adapter_050:source0_endofpacket -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_050_source0_valid;                                                         // burst_adapter_050:source0_valid -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_050_source0_startofpacket;                                                 // burst_adapter_050:source0_startofpacket -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_050_source0_data;                                                          // burst_adapter_050:source0_data -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_050_source0_ready;                                                         // Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_050:source0_ready
	wire  [57:0] burst_adapter_050_source0_channel;                                                       // burst_adapter_050:source0_channel -> Shiled_IO_A23_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         burst_adapter_051_source0_endofpacket;                                                   // burst_adapter_051:source0_endofpacket -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_051_source0_valid;                                                         // burst_adapter_051:source0_valid -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_051_source0_startofpacket;                                                 // burst_adapter_051:source0_startofpacket -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [65:0] burst_adapter_051_source0_data;                                                          // burst_adapter_051:source0_data -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_051_source0_ready;                                                         // Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_051:source0_ready
	wire  [57:0] burst_adapter_051_source0_channel;                                                       // burst_adapter_051:source0_channel -> Shiled_IO_A18_ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src0_endofpacket;                                                         // cmd_xbar_demux:src0_endofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                               // cmd_xbar_demux:src0_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                       // cmd_xbar_demux:src0_startofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_src0_data;                                                                // cmd_xbar_demux:src0_data -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_data
	wire  [57:0] cmd_xbar_demux_src0_channel;                                                             // cmd_xbar_demux:src0_channel -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src1_endofpacket;                                                         // cmd_xbar_demux:src1_endofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                               // cmd_xbar_demux:src1_valid -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                       // cmd_xbar_demux:src1_startofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_src1_data;                                                                // cmd_xbar_demux:src1_data -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire  [57:0] cmd_xbar_demux_src1_channel;                                                             // cmd_xbar_demux:src1_channel -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src2_endofpacket;                                                         // cmd_xbar_demux:src2_endofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                               // cmd_xbar_demux:src2_valid -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                       // cmd_xbar_demux:src2_startofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_src2_data;                                                                // cmd_xbar_demux:src2_data -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire  [57:0] cmd_xbar_demux_src2_channel;                                                             // cmd_xbar_demux:src2_channel -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src3_endofpacket;                                                         // cmd_xbar_demux:src3_endofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                               // cmd_xbar_demux:src3_valid -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                       // cmd_xbar_demux:src3_startofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_src3_data;                                                                // cmd_xbar_demux:src3_data -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire  [57:0] cmd_xbar_demux_src3_channel;                                                             // cmd_xbar_demux:src3_channel -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src4_endofpacket;                                                         // cmd_xbar_demux:src4_endofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                               // cmd_xbar_demux:src4_valid -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                       // cmd_xbar_demux:src4_startofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_src4_data;                                                                // cmd_xbar_demux:src4_data -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire  [57:0] cmd_xbar_demux_src4_channel;                                                             // cmd_xbar_demux:src4_channel -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src5_endofpacket;                                                         // cmd_xbar_demux:src5_endofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src5_valid;                                                               // cmd_xbar_demux:src5_valid -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src5_startofpacket;                                                       // cmd_xbar_demux:src5_startofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_demux_src5_data;                                                                // cmd_xbar_demux:src5_data -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire  [57:0] cmd_xbar_demux_src5_channel;                                                             // cmd_xbar_demux:src5_channel -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src6_endofpacket;                                                         // cmd_xbar_demux:src6_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_demux_src6_valid;                                                               // cmd_xbar_demux:src6_valid -> width_adapter:in_valid
	wire         cmd_xbar_demux_src6_startofpacket;                                                       // cmd_xbar_demux:src6_startofpacket -> width_adapter:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src6_data;                                                                // cmd_xbar_demux:src6_data -> width_adapter:in_data
	wire  [57:0] cmd_xbar_demux_src6_channel;                                                             // cmd_xbar_demux:src6_channel -> width_adapter:in_channel
	wire         cmd_xbar_demux_src7_endofpacket;                                                         // cmd_xbar_demux:src7_endofpacket -> width_adapter_002:in_endofpacket
	wire         cmd_xbar_demux_src7_valid;                                                               // cmd_xbar_demux:src7_valid -> width_adapter_002:in_valid
	wire         cmd_xbar_demux_src7_startofpacket;                                                       // cmd_xbar_demux:src7_startofpacket -> width_adapter_002:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src7_data;                                                                // cmd_xbar_demux:src7_data -> width_adapter_002:in_data
	wire  [57:0] cmd_xbar_demux_src7_channel;                                                             // cmd_xbar_demux:src7_channel -> width_adapter_002:in_channel
	wire         cmd_xbar_demux_src8_endofpacket;                                                         // cmd_xbar_demux:src8_endofpacket -> width_adapter_004:in_endofpacket
	wire         cmd_xbar_demux_src8_valid;                                                               // cmd_xbar_demux:src8_valid -> width_adapter_004:in_valid
	wire         cmd_xbar_demux_src8_startofpacket;                                                       // cmd_xbar_demux:src8_startofpacket -> width_adapter_004:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src8_data;                                                                // cmd_xbar_demux:src8_data -> width_adapter_004:in_data
	wire  [57:0] cmd_xbar_demux_src8_channel;                                                             // cmd_xbar_demux:src8_channel -> width_adapter_004:in_channel
	wire         cmd_xbar_demux_src9_endofpacket;                                                         // cmd_xbar_demux:src9_endofpacket -> width_adapter_006:in_endofpacket
	wire         cmd_xbar_demux_src9_valid;                                                               // cmd_xbar_demux:src9_valid -> width_adapter_006:in_valid
	wire         cmd_xbar_demux_src9_startofpacket;                                                       // cmd_xbar_demux:src9_startofpacket -> width_adapter_006:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src9_data;                                                                // cmd_xbar_demux:src9_data -> width_adapter_006:in_data
	wire  [57:0] cmd_xbar_demux_src9_channel;                                                             // cmd_xbar_demux:src9_channel -> width_adapter_006:in_channel
	wire         cmd_xbar_demux_src10_endofpacket;                                                        // cmd_xbar_demux:src10_endofpacket -> width_adapter_008:in_endofpacket
	wire         cmd_xbar_demux_src10_valid;                                                              // cmd_xbar_demux:src10_valid -> width_adapter_008:in_valid
	wire         cmd_xbar_demux_src10_startofpacket;                                                      // cmd_xbar_demux:src10_startofpacket -> width_adapter_008:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src10_data;                                                               // cmd_xbar_demux:src10_data -> width_adapter_008:in_data
	wire  [57:0] cmd_xbar_demux_src10_channel;                                                            // cmd_xbar_demux:src10_channel -> width_adapter_008:in_channel
	wire         cmd_xbar_demux_src11_endofpacket;                                                        // cmd_xbar_demux:src11_endofpacket -> width_adapter_010:in_endofpacket
	wire         cmd_xbar_demux_src11_valid;                                                              // cmd_xbar_demux:src11_valid -> width_adapter_010:in_valid
	wire         cmd_xbar_demux_src11_startofpacket;                                                      // cmd_xbar_demux:src11_startofpacket -> width_adapter_010:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src11_data;                                                               // cmd_xbar_demux:src11_data -> width_adapter_010:in_data
	wire  [57:0] cmd_xbar_demux_src11_channel;                                                            // cmd_xbar_demux:src11_channel -> width_adapter_010:in_channel
	wire         cmd_xbar_demux_src12_endofpacket;                                                        // cmd_xbar_demux:src12_endofpacket -> width_adapter_012:in_endofpacket
	wire         cmd_xbar_demux_src12_valid;                                                              // cmd_xbar_demux:src12_valid -> width_adapter_012:in_valid
	wire         cmd_xbar_demux_src12_startofpacket;                                                      // cmd_xbar_demux:src12_startofpacket -> width_adapter_012:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src12_data;                                                               // cmd_xbar_demux:src12_data -> width_adapter_012:in_data
	wire  [57:0] cmd_xbar_demux_src12_channel;                                                            // cmd_xbar_demux:src12_channel -> width_adapter_012:in_channel
	wire         cmd_xbar_demux_src13_endofpacket;                                                        // cmd_xbar_demux:src13_endofpacket -> width_adapter_014:in_endofpacket
	wire         cmd_xbar_demux_src13_valid;                                                              // cmd_xbar_demux:src13_valid -> width_adapter_014:in_valid
	wire         cmd_xbar_demux_src13_startofpacket;                                                      // cmd_xbar_demux:src13_startofpacket -> width_adapter_014:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src13_data;                                                               // cmd_xbar_demux:src13_data -> width_adapter_014:in_data
	wire  [57:0] cmd_xbar_demux_src13_channel;                                                            // cmd_xbar_demux:src13_channel -> width_adapter_014:in_channel
	wire         cmd_xbar_demux_src14_endofpacket;                                                        // cmd_xbar_demux:src14_endofpacket -> width_adapter_016:in_endofpacket
	wire         cmd_xbar_demux_src14_valid;                                                              // cmd_xbar_demux:src14_valid -> width_adapter_016:in_valid
	wire         cmd_xbar_demux_src14_startofpacket;                                                      // cmd_xbar_demux:src14_startofpacket -> width_adapter_016:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src14_data;                                                               // cmd_xbar_demux:src14_data -> width_adapter_016:in_data
	wire  [57:0] cmd_xbar_demux_src14_channel;                                                            // cmd_xbar_demux:src14_channel -> width_adapter_016:in_channel
	wire         cmd_xbar_demux_src15_endofpacket;                                                        // cmd_xbar_demux:src15_endofpacket -> width_adapter_018:in_endofpacket
	wire         cmd_xbar_demux_src15_valid;                                                              // cmd_xbar_demux:src15_valid -> width_adapter_018:in_valid
	wire         cmd_xbar_demux_src15_startofpacket;                                                      // cmd_xbar_demux:src15_startofpacket -> width_adapter_018:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src15_data;                                                               // cmd_xbar_demux:src15_data -> width_adapter_018:in_data
	wire  [57:0] cmd_xbar_demux_src15_channel;                                                            // cmd_xbar_demux:src15_channel -> width_adapter_018:in_channel
	wire         cmd_xbar_demux_src16_endofpacket;                                                        // cmd_xbar_demux:src16_endofpacket -> width_adapter_020:in_endofpacket
	wire         cmd_xbar_demux_src16_valid;                                                              // cmd_xbar_demux:src16_valid -> width_adapter_020:in_valid
	wire         cmd_xbar_demux_src16_startofpacket;                                                      // cmd_xbar_demux:src16_startofpacket -> width_adapter_020:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src16_data;                                                               // cmd_xbar_demux:src16_data -> width_adapter_020:in_data
	wire  [57:0] cmd_xbar_demux_src16_channel;                                                            // cmd_xbar_demux:src16_channel -> width_adapter_020:in_channel
	wire         cmd_xbar_demux_src17_endofpacket;                                                        // cmd_xbar_demux:src17_endofpacket -> width_adapter_022:in_endofpacket
	wire         cmd_xbar_demux_src17_valid;                                                              // cmd_xbar_demux:src17_valid -> width_adapter_022:in_valid
	wire         cmd_xbar_demux_src17_startofpacket;                                                      // cmd_xbar_demux:src17_startofpacket -> width_adapter_022:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src17_data;                                                               // cmd_xbar_demux:src17_data -> width_adapter_022:in_data
	wire  [57:0] cmd_xbar_demux_src17_channel;                                                            // cmd_xbar_demux:src17_channel -> width_adapter_022:in_channel
	wire         cmd_xbar_demux_src18_endofpacket;                                                        // cmd_xbar_demux:src18_endofpacket -> width_adapter_024:in_endofpacket
	wire         cmd_xbar_demux_src18_valid;                                                              // cmd_xbar_demux:src18_valid -> width_adapter_024:in_valid
	wire         cmd_xbar_demux_src18_startofpacket;                                                      // cmd_xbar_demux:src18_startofpacket -> width_adapter_024:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src18_data;                                                               // cmd_xbar_demux:src18_data -> width_adapter_024:in_data
	wire  [57:0] cmd_xbar_demux_src18_channel;                                                            // cmd_xbar_demux:src18_channel -> width_adapter_024:in_channel
	wire         cmd_xbar_demux_src19_endofpacket;                                                        // cmd_xbar_demux:src19_endofpacket -> width_adapter_026:in_endofpacket
	wire         cmd_xbar_demux_src19_valid;                                                              // cmd_xbar_demux:src19_valid -> width_adapter_026:in_valid
	wire         cmd_xbar_demux_src19_startofpacket;                                                      // cmd_xbar_demux:src19_startofpacket -> width_adapter_026:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src19_data;                                                               // cmd_xbar_demux:src19_data -> width_adapter_026:in_data
	wire  [57:0] cmd_xbar_demux_src19_channel;                                                            // cmd_xbar_demux:src19_channel -> width_adapter_026:in_channel
	wire         cmd_xbar_demux_src20_endofpacket;                                                        // cmd_xbar_demux:src20_endofpacket -> width_adapter_028:in_endofpacket
	wire         cmd_xbar_demux_src20_valid;                                                              // cmd_xbar_demux:src20_valid -> width_adapter_028:in_valid
	wire         cmd_xbar_demux_src20_startofpacket;                                                      // cmd_xbar_demux:src20_startofpacket -> width_adapter_028:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src20_data;                                                               // cmd_xbar_demux:src20_data -> width_adapter_028:in_data
	wire  [57:0] cmd_xbar_demux_src20_channel;                                                            // cmd_xbar_demux:src20_channel -> width_adapter_028:in_channel
	wire         cmd_xbar_demux_src21_endofpacket;                                                        // cmd_xbar_demux:src21_endofpacket -> width_adapter_030:in_endofpacket
	wire         cmd_xbar_demux_src21_valid;                                                              // cmd_xbar_demux:src21_valid -> width_adapter_030:in_valid
	wire         cmd_xbar_demux_src21_startofpacket;                                                      // cmd_xbar_demux:src21_startofpacket -> width_adapter_030:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src21_data;                                                               // cmd_xbar_demux:src21_data -> width_adapter_030:in_data
	wire  [57:0] cmd_xbar_demux_src21_channel;                                                            // cmd_xbar_demux:src21_channel -> width_adapter_030:in_channel
	wire         cmd_xbar_demux_src22_endofpacket;                                                        // cmd_xbar_demux:src22_endofpacket -> width_adapter_032:in_endofpacket
	wire         cmd_xbar_demux_src22_valid;                                                              // cmd_xbar_demux:src22_valid -> width_adapter_032:in_valid
	wire         cmd_xbar_demux_src22_startofpacket;                                                      // cmd_xbar_demux:src22_startofpacket -> width_adapter_032:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src22_data;                                                               // cmd_xbar_demux:src22_data -> width_adapter_032:in_data
	wire  [57:0] cmd_xbar_demux_src22_channel;                                                            // cmd_xbar_demux:src22_channel -> width_adapter_032:in_channel
	wire         cmd_xbar_demux_src23_endofpacket;                                                        // cmd_xbar_demux:src23_endofpacket -> width_adapter_034:in_endofpacket
	wire         cmd_xbar_demux_src23_valid;                                                              // cmd_xbar_demux:src23_valid -> width_adapter_034:in_valid
	wire         cmd_xbar_demux_src23_startofpacket;                                                      // cmd_xbar_demux:src23_startofpacket -> width_adapter_034:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src23_data;                                                               // cmd_xbar_demux:src23_data -> width_adapter_034:in_data
	wire  [57:0] cmd_xbar_demux_src23_channel;                                                            // cmd_xbar_demux:src23_channel -> width_adapter_034:in_channel
	wire         cmd_xbar_demux_src24_endofpacket;                                                        // cmd_xbar_demux:src24_endofpacket -> width_adapter_036:in_endofpacket
	wire         cmd_xbar_demux_src24_valid;                                                              // cmd_xbar_demux:src24_valid -> width_adapter_036:in_valid
	wire         cmd_xbar_demux_src24_startofpacket;                                                      // cmd_xbar_demux:src24_startofpacket -> width_adapter_036:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src24_data;                                                               // cmd_xbar_demux:src24_data -> width_adapter_036:in_data
	wire  [57:0] cmd_xbar_demux_src24_channel;                                                            // cmd_xbar_demux:src24_channel -> width_adapter_036:in_channel
	wire         cmd_xbar_demux_src25_endofpacket;                                                        // cmd_xbar_demux:src25_endofpacket -> width_adapter_038:in_endofpacket
	wire         cmd_xbar_demux_src25_valid;                                                              // cmd_xbar_demux:src25_valid -> width_adapter_038:in_valid
	wire         cmd_xbar_demux_src25_startofpacket;                                                      // cmd_xbar_demux:src25_startofpacket -> width_adapter_038:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src25_data;                                                               // cmd_xbar_demux:src25_data -> width_adapter_038:in_data
	wire  [57:0] cmd_xbar_demux_src25_channel;                                                            // cmd_xbar_demux:src25_channel -> width_adapter_038:in_channel
	wire         cmd_xbar_demux_src26_endofpacket;                                                        // cmd_xbar_demux:src26_endofpacket -> width_adapter_040:in_endofpacket
	wire         cmd_xbar_demux_src26_valid;                                                              // cmd_xbar_demux:src26_valid -> width_adapter_040:in_valid
	wire         cmd_xbar_demux_src26_startofpacket;                                                      // cmd_xbar_demux:src26_startofpacket -> width_adapter_040:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src26_data;                                                               // cmd_xbar_demux:src26_data -> width_adapter_040:in_data
	wire  [57:0] cmd_xbar_demux_src26_channel;                                                            // cmd_xbar_demux:src26_channel -> width_adapter_040:in_channel
	wire         cmd_xbar_demux_src27_endofpacket;                                                        // cmd_xbar_demux:src27_endofpacket -> width_adapter_042:in_endofpacket
	wire         cmd_xbar_demux_src27_valid;                                                              // cmd_xbar_demux:src27_valid -> width_adapter_042:in_valid
	wire         cmd_xbar_demux_src27_startofpacket;                                                      // cmd_xbar_demux:src27_startofpacket -> width_adapter_042:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src27_data;                                                               // cmd_xbar_demux:src27_data -> width_adapter_042:in_data
	wire  [57:0] cmd_xbar_demux_src27_channel;                                                            // cmd_xbar_demux:src27_channel -> width_adapter_042:in_channel
	wire         cmd_xbar_demux_src28_endofpacket;                                                        // cmd_xbar_demux:src28_endofpacket -> width_adapter_044:in_endofpacket
	wire         cmd_xbar_demux_src28_valid;                                                              // cmd_xbar_demux:src28_valid -> width_adapter_044:in_valid
	wire         cmd_xbar_demux_src28_startofpacket;                                                      // cmd_xbar_demux:src28_startofpacket -> width_adapter_044:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src28_data;                                                               // cmd_xbar_demux:src28_data -> width_adapter_044:in_data
	wire  [57:0] cmd_xbar_demux_src28_channel;                                                            // cmd_xbar_demux:src28_channel -> width_adapter_044:in_channel
	wire         cmd_xbar_demux_src29_endofpacket;                                                        // cmd_xbar_demux:src29_endofpacket -> width_adapter_046:in_endofpacket
	wire         cmd_xbar_demux_src29_valid;                                                              // cmd_xbar_demux:src29_valid -> width_adapter_046:in_valid
	wire         cmd_xbar_demux_src29_startofpacket;                                                      // cmd_xbar_demux:src29_startofpacket -> width_adapter_046:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src29_data;                                                               // cmd_xbar_demux:src29_data -> width_adapter_046:in_data
	wire  [57:0] cmd_xbar_demux_src29_channel;                                                            // cmd_xbar_demux:src29_channel -> width_adapter_046:in_channel
	wire         cmd_xbar_demux_src30_endofpacket;                                                        // cmd_xbar_demux:src30_endofpacket -> width_adapter_048:in_endofpacket
	wire         cmd_xbar_demux_src30_valid;                                                              // cmd_xbar_demux:src30_valid -> width_adapter_048:in_valid
	wire         cmd_xbar_demux_src30_startofpacket;                                                      // cmd_xbar_demux:src30_startofpacket -> width_adapter_048:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src30_data;                                                               // cmd_xbar_demux:src30_data -> width_adapter_048:in_data
	wire  [57:0] cmd_xbar_demux_src30_channel;                                                            // cmd_xbar_demux:src30_channel -> width_adapter_048:in_channel
	wire         cmd_xbar_demux_src31_endofpacket;                                                        // cmd_xbar_demux:src31_endofpacket -> width_adapter_050:in_endofpacket
	wire         cmd_xbar_demux_src31_valid;                                                              // cmd_xbar_demux:src31_valid -> width_adapter_050:in_valid
	wire         cmd_xbar_demux_src31_startofpacket;                                                      // cmd_xbar_demux:src31_startofpacket -> width_adapter_050:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src31_data;                                                               // cmd_xbar_demux:src31_data -> width_adapter_050:in_data
	wire  [57:0] cmd_xbar_demux_src31_channel;                                                            // cmd_xbar_demux:src31_channel -> width_adapter_050:in_channel
	wire         cmd_xbar_demux_src32_endofpacket;                                                        // cmd_xbar_demux:src32_endofpacket -> width_adapter_052:in_endofpacket
	wire         cmd_xbar_demux_src32_valid;                                                              // cmd_xbar_demux:src32_valid -> width_adapter_052:in_valid
	wire         cmd_xbar_demux_src32_startofpacket;                                                      // cmd_xbar_demux:src32_startofpacket -> width_adapter_052:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src32_data;                                                               // cmd_xbar_demux:src32_data -> width_adapter_052:in_data
	wire  [57:0] cmd_xbar_demux_src32_channel;                                                            // cmd_xbar_demux:src32_channel -> width_adapter_052:in_channel
	wire         cmd_xbar_demux_src33_endofpacket;                                                        // cmd_xbar_demux:src33_endofpacket -> width_adapter_054:in_endofpacket
	wire         cmd_xbar_demux_src33_valid;                                                              // cmd_xbar_demux:src33_valid -> width_adapter_054:in_valid
	wire         cmd_xbar_demux_src33_startofpacket;                                                      // cmd_xbar_demux:src33_startofpacket -> width_adapter_054:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src33_data;                                                               // cmd_xbar_demux:src33_data -> width_adapter_054:in_data
	wire  [57:0] cmd_xbar_demux_src33_channel;                                                            // cmd_xbar_demux:src33_channel -> width_adapter_054:in_channel
	wire         cmd_xbar_demux_src34_endofpacket;                                                        // cmd_xbar_demux:src34_endofpacket -> width_adapter_056:in_endofpacket
	wire         cmd_xbar_demux_src34_valid;                                                              // cmd_xbar_demux:src34_valid -> width_adapter_056:in_valid
	wire         cmd_xbar_demux_src34_startofpacket;                                                      // cmd_xbar_demux:src34_startofpacket -> width_adapter_056:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src34_data;                                                               // cmd_xbar_demux:src34_data -> width_adapter_056:in_data
	wire  [57:0] cmd_xbar_demux_src34_channel;                                                            // cmd_xbar_demux:src34_channel -> width_adapter_056:in_channel
	wire         cmd_xbar_demux_src35_endofpacket;                                                        // cmd_xbar_demux:src35_endofpacket -> width_adapter_058:in_endofpacket
	wire         cmd_xbar_demux_src35_valid;                                                              // cmd_xbar_demux:src35_valid -> width_adapter_058:in_valid
	wire         cmd_xbar_demux_src35_startofpacket;                                                      // cmd_xbar_demux:src35_startofpacket -> width_adapter_058:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src35_data;                                                               // cmd_xbar_demux:src35_data -> width_adapter_058:in_data
	wire  [57:0] cmd_xbar_demux_src35_channel;                                                            // cmd_xbar_demux:src35_channel -> width_adapter_058:in_channel
	wire         cmd_xbar_demux_src36_endofpacket;                                                        // cmd_xbar_demux:src36_endofpacket -> width_adapter_060:in_endofpacket
	wire         cmd_xbar_demux_src36_valid;                                                              // cmd_xbar_demux:src36_valid -> width_adapter_060:in_valid
	wire         cmd_xbar_demux_src36_startofpacket;                                                      // cmd_xbar_demux:src36_startofpacket -> width_adapter_060:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src36_data;                                                               // cmd_xbar_demux:src36_data -> width_adapter_060:in_data
	wire  [57:0] cmd_xbar_demux_src36_channel;                                                            // cmd_xbar_demux:src36_channel -> width_adapter_060:in_channel
	wire         cmd_xbar_demux_src37_endofpacket;                                                        // cmd_xbar_demux:src37_endofpacket -> width_adapter_062:in_endofpacket
	wire         cmd_xbar_demux_src37_valid;                                                              // cmd_xbar_demux:src37_valid -> width_adapter_062:in_valid
	wire         cmd_xbar_demux_src37_startofpacket;                                                      // cmd_xbar_demux:src37_startofpacket -> width_adapter_062:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src37_data;                                                               // cmd_xbar_demux:src37_data -> width_adapter_062:in_data
	wire  [57:0] cmd_xbar_demux_src37_channel;                                                            // cmd_xbar_demux:src37_channel -> width_adapter_062:in_channel
	wire         cmd_xbar_demux_src38_endofpacket;                                                        // cmd_xbar_demux:src38_endofpacket -> width_adapter_064:in_endofpacket
	wire         cmd_xbar_demux_src38_valid;                                                              // cmd_xbar_demux:src38_valid -> width_adapter_064:in_valid
	wire         cmd_xbar_demux_src38_startofpacket;                                                      // cmd_xbar_demux:src38_startofpacket -> width_adapter_064:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src38_data;                                                               // cmd_xbar_demux:src38_data -> width_adapter_064:in_data
	wire  [57:0] cmd_xbar_demux_src38_channel;                                                            // cmd_xbar_demux:src38_channel -> width_adapter_064:in_channel
	wire         cmd_xbar_demux_src39_endofpacket;                                                        // cmd_xbar_demux:src39_endofpacket -> width_adapter_066:in_endofpacket
	wire         cmd_xbar_demux_src39_valid;                                                              // cmd_xbar_demux:src39_valid -> width_adapter_066:in_valid
	wire         cmd_xbar_demux_src39_startofpacket;                                                      // cmd_xbar_demux:src39_startofpacket -> width_adapter_066:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src39_data;                                                               // cmd_xbar_demux:src39_data -> width_adapter_066:in_data
	wire  [57:0] cmd_xbar_demux_src39_channel;                                                            // cmd_xbar_demux:src39_channel -> width_adapter_066:in_channel
	wire         cmd_xbar_demux_src40_endofpacket;                                                        // cmd_xbar_demux:src40_endofpacket -> width_adapter_068:in_endofpacket
	wire         cmd_xbar_demux_src40_valid;                                                              // cmd_xbar_demux:src40_valid -> width_adapter_068:in_valid
	wire         cmd_xbar_demux_src40_startofpacket;                                                      // cmd_xbar_demux:src40_startofpacket -> width_adapter_068:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src40_data;                                                               // cmd_xbar_demux:src40_data -> width_adapter_068:in_data
	wire  [57:0] cmd_xbar_demux_src40_channel;                                                            // cmd_xbar_demux:src40_channel -> width_adapter_068:in_channel
	wire         cmd_xbar_demux_src41_endofpacket;                                                        // cmd_xbar_demux:src41_endofpacket -> width_adapter_070:in_endofpacket
	wire         cmd_xbar_demux_src41_valid;                                                              // cmd_xbar_demux:src41_valid -> width_adapter_070:in_valid
	wire         cmd_xbar_demux_src41_startofpacket;                                                      // cmd_xbar_demux:src41_startofpacket -> width_adapter_070:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src41_data;                                                               // cmd_xbar_demux:src41_data -> width_adapter_070:in_data
	wire  [57:0] cmd_xbar_demux_src41_channel;                                                            // cmd_xbar_demux:src41_channel -> width_adapter_070:in_channel
	wire         cmd_xbar_demux_src42_endofpacket;                                                        // cmd_xbar_demux:src42_endofpacket -> width_adapter_072:in_endofpacket
	wire         cmd_xbar_demux_src42_valid;                                                              // cmd_xbar_demux:src42_valid -> width_adapter_072:in_valid
	wire         cmd_xbar_demux_src42_startofpacket;                                                      // cmd_xbar_demux:src42_startofpacket -> width_adapter_072:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src42_data;                                                               // cmd_xbar_demux:src42_data -> width_adapter_072:in_data
	wire  [57:0] cmd_xbar_demux_src42_channel;                                                            // cmd_xbar_demux:src42_channel -> width_adapter_072:in_channel
	wire         cmd_xbar_demux_src43_endofpacket;                                                        // cmd_xbar_demux:src43_endofpacket -> width_adapter_074:in_endofpacket
	wire         cmd_xbar_demux_src43_valid;                                                              // cmd_xbar_demux:src43_valid -> width_adapter_074:in_valid
	wire         cmd_xbar_demux_src43_startofpacket;                                                      // cmd_xbar_demux:src43_startofpacket -> width_adapter_074:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src43_data;                                                               // cmd_xbar_demux:src43_data -> width_adapter_074:in_data
	wire  [57:0] cmd_xbar_demux_src43_channel;                                                            // cmd_xbar_demux:src43_channel -> width_adapter_074:in_channel
	wire         cmd_xbar_demux_src44_endofpacket;                                                        // cmd_xbar_demux:src44_endofpacket -> width_adapter_076:in_endofpacket
	wire         cmd_xbar_demux_src44_valid;                                                              // cmd_xbar_demux:src44_valid -> width_adapter_076:in_valid
	wire         cmd_xbar_demux_src44_startofpacket;                                                      // cmd_xbar_demux:src44_startofpacket -> width_adapter_076:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src44_data;                                                               // cmd_xbar_demux:src44_data -> width_adapter_076:in_data
	wire  [57:0] cmd_xbar_demux_src44_channel;                                                            // cmd_xbar_demux:src44_channel -> width_adapter_076:in_channel
	wire         cmd_xbar_demux_src45_endofpacket;                                                        // cmd_xbar_demux:src45_endofpacket -> width_adapter_078:in_endofpacket
	wire         cmd_xbar_demux_src45_valid;                                                              // cmd_xbar_demux:src45_valid -> width_adapter_078:in_valid
	wire         cmd_xbar_demux_src45_startofpacket;                                                      // cmd_xbar_demux:src45_startofpacket -> width_adapter_078:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src45_data;                                                               // cmd_xbar_demux:src45_data -> width_adapter_078:in_data
	wire  [57:0] cmd_xbar_demux_src45_channel;                                                            // cmd_xbar_demux:src45_channel -> width_adapter_078:in_channel
	wire         cmd_xbar_demux_src46_endofpacket;                                                        // cmd_xbar_demux:src46_endofpacket -> width_adapter_080:in_endofpacket
	wire         cmd_xbar_demux_src46_valid;                                                              // cmd_xbar_demux:src46_valid -> width_adapter_080:in_valid
	wire         cmd_xbar_demux_src46_startofpacket;                                                      // cmd_xbar_demux:src46_startofpacket -> width_adapter_080:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src46_data;                                                               // cmd_xbar_demux:src46_data -> width_adapter_080:in_data
	wire  [57:0] cmd_xbar_demux_src46_channel;                                                            // cmd_xbar_demux:src46_channel -> width_adapter_080:in_channel
	wire         cmd_xbar_demux_src47_endofpacket;                                                        // cmd_xbar_demux:src47_endofpacket -> width_adapter_082:in_endofpacket
	wire         cmd_xbar_demux_src47_valid;                                                              // cmd_xbar_demux:src47_valid -> width_adapter_082:in_valid
	wire         cmd_xbar_demux_src47_startofpacket;                                                      // cmd_xbar_demux:src47_startofpacket -> width_adapter_082:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src47_data;                                                               // cmd_xbar_demux:src47_data -> width_adapter_082:in_data
	wire  [57:0] cmd_xbar_demux_src47_channel;                                                            // cmd_xbar_demux:src47_channel -> width_adapter_082:in_channel
	wire         cmd_xbar_demux_src48_endofpacket;                                                        // cmd_xbar_demux:src48_endofpacket -> width_adapter_084:in_endofpacket
	wire         cmd_xbar_demux_src48_valid;                                                              // cmd_xbar_demux:src48_valid -> width_adapter_084:in_valid
	wire         cmd_xbar_demux_src48_startofpacket;                                                      // cmd_xbar_demux:src48_startofpacket -> width_adapter_084:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src48_data;                                                               // cmd_xbar_demux:src48_data -> width_adapter_084:in_data
	wire  [57:0] cmd_xbar_demux_src48_channel;                                                            // cmd_xbar_demux:src48_channel -> width_adapter_084:in_channel
	wire         cmd_xbar_demux_src49_endofpacket;                                                        // cmd_xbar_demux:src49_endofpacket -> width_adapter_086:in_endofpacket
	wire         cmd_xbar_demux_src49_valid;                                                              // cmd_xbar_demux:src49_valid -> width_adapter_086:in_valid
	wire         cmd_xbar_demux_src49_startofpacket;                                                      // cmd_xbar_demux:src49_startofpacket -> width_adapter_086:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src49_data;                                                               // cmd_xbar_demux:src49_data -> width_adapter_086:in_data
	wire  [57:0] cmd_xbar_demux_src49_channel;                                                            // cmd_xbar_demux:src49_channel -> width_adapter_086:in_channel
	wire         cmd_xbar_demux_src50_endofpacket;                                                        // cmd_xbar_demux:src50_endofpacket -> width_adapter_088:in_endofpacket
	wire         cmd_xbar_demux_src50_valid;                                                              // cmd_xbar_demux:src50_valid -> width_adapter_088:in_valid
	wire         cmd_xbar_demux_src50_startofpacket;                                                      // cmd_xbar_demux:src50_startofpacket -> width_adapter_088:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src50_data;                                                               // cmd_xbar_demux:src50_data -> width_adapter_088:in_data
	wire  [57:0] cmd_xbar_demux_src50_channel;                                                            // cmd_xbar_demux:src50_channel -> width_adapter_088:in_channel
	wire         cmd_xbar_demux_src51_endofpacket;                                                        // cmd_xbar_demux:src51_endofpacket -> width_adapter_090:in_endofpacket
	wire         cmd_xbar_demux_src51_valid;                                                              // cmd_xbar_demux:src51_valid -> width_adapter_090:in_valid
	wire         cmd_xbar_demux_src51_startofpacket;                                                      // cmd_xbar_demux:src51_startofpacket -> width_adapter_090:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src51_data;                                                               // cmd_xbar_demux:src51_data -> width_adapter_090:in_data
	wire  [57:0] cmd_xbar_demux_src51_channel;                                                            // cmd_xbar_demux:src51_channel -> width_adapter_090:in_channel
	wire         cmd_xbar_demux_src52_endofpacket;                                                        // cmd_xbar_demux:src52_endofpacket -> width_adapter_092:in_endofpacket
	wire         cmd_xbar_demux_src52_valid;                                                              // cmd_xbar_demux:src52_valid -> width_adapter_092:in_valid
	wire         cmd_xbar_demux_src52_startofpacket;                                                      // cmd_xbar_demux:src52_startofpacket -> width_adapter_092:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src52_data;                                                               // cmd_xbar_demux:src52_data -> width_adapter_092:in_data
	wire  [57:0] cmd_xbar_demux_src52_channel;                                                            // cmd_xbar_demux:src52_channel -> width_adapter_092:in_channel
	wire         cmd_xbar_demux_src53_endofpacket;                                                        // cmd_xbar_demux:src53_endofpacket -> width_adapter_094:in_endofpacket
	wire         cmd_xbar_demux_src53_valid;                                                              // cmd_xbar_demux:src53_valid -> width_adapter_094:in_valid
	wire         cmd_xbar_demux_src53_startofpacket;                                                      // cmd_xbar_demux:src53_startofpacket -> width_adapter_094:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src53_data;                                                               // cmd_xbar_demux:src53_data -> width_adapter_094:in_data
	wire  [57:0] cmd_xbar_demux_src53_channel;                                                            // cmd_xbar_demux:src53_channel -> width_adapter_094:in_channel
	wire         cmd_xbar_demux_src54_endofpacket;                                                        // cmd_xbar_demux:src54_endofpacket -> width_adapter_096:in_endofpacket
	wire         cmd_xbar_demux_src54_valid;                                                              // cmd_xbar_demux:src54_valid -> width_adapter_096:in_valid
	wire         cmd_xbar_demux_src54_startofpacket;                                                      // cmd_xbar_demux:src54_startofpacket -> width_adapter_096:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src54_data;                                                               // cmd_xbar_demux:src54_data -> width_adapter_096:in_data
	wire  [57:0] cmd_xbar_demux_src54_channel;                                                            // cmd_xbar_demux:src54_channel -> width_adapter_096:in_channel
	wire         cmd_xbar_demux_src55_endofpacket;                                                        // cmd_xbar_demux:src55_endofpacket -> width_adapter_098:in_endofpacket
	wire         cmd_xbar_demux_src55_valid;                                                              // cmd_xbar_demux:src55_valid -> width_adapter_098:in_valid
	wire         cmd_xbar_demux_src55_startofpacket;                                                      // cmd_xbar_demux:src55_startofpacket -> width_adapter_098:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src55_data;                                                               // cmd_xbar_demux:src55_data -> width_adapter_098:in_data
	wire  [57:0] cmd_xbar_demux_src55_channel;                                                            // cmd_xbar_demux:src55_channel -> width_adapter_098:in_channel
	wire         cmd_xbar_demux_src56_endofpacket;                                                        // cmd_xbar_demux:src56_endofpacket -> width_adapter_100:in_endofpacket
	wire         cmd_xbar_demux_src56_valid;                                                              // cmd_xbar_demux:src56_valid -> width_adapter_100:in_valid
	wire         cmd_xbar_demux_src56_startofpacket;                                                      // cmd_xbar_demux:src56_startofpacket -> width_adapter_100:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src56_data;                                                               // cmd_xbar_demux:src56_data -> width_adapter_100:in_data
	wire  [57:0] cmd_xbar_demux_src56_channel;                                                            // cmd_xbar_demux:src56_channel -> width_adapter_100:in_channel
	wire         cmd_xbar_demux_src57_endofpacket;                                                        // cmd_xbar_demux:src57_endofpacket -> width_adapter_102:in_endofpacket
	wire         cmd_xbar_demux_src57_valid;                                                              // cmd_xbar_demux:src57_valid -> width_adapter_102:in_valid
	wire         cmd_xbar_demux_src57_startofpacket;                                                      // cmd_xbar_demux:src57_startofpacket -> width_adapter_102:in_startofpacket
	wire  [92:0] cmd_xbar_demux_src57_data;                                                               // cmd_xbar_demux:src57_data -> width_adapter_102:in_data
	wire  [57:0] cmd_xbar_demux_src57_channel;                                                            // cmd_xbar_demux:src57_channel -> width_adapter_102:in_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                         // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                               // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                       // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [92:0] rsp_xbar_demux_src0_data;                                                                // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [57:0] rsp_xbar_demux_src0_channel;                                                             // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                               // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                     // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                           // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                   // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [92:0] rsp_xbar_demux_001_src0_data;                                                            // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [57:0] rsp_xbar_demux_001_src0_channel;                                                         // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                           // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                     // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                           // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                   // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [92:0] rsp_xbar_demux_002_src0_data;                                                            // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [57:0] rsp_xbar_demux_002_src0_channel;                                                         // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                           // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                     // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                           // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                   // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [92:0] rsp_xbar_demux_003_src0_data;                                                            // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire  [57:0] rsp_xbar_demux_003_src0_channel;                                                         // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                           // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                     // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                           // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                   // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [92:0] rsp_xbar_demux_004_src0_data;                                                            // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire  [57:0] rsp_xbar_demux_004_src0_channel;                                                         // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                           // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                     // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                           // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                   // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [92:0] rsp_xbar_demux_005_src0_data;                                                            // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire  [57:0] rsp_xbar_demux_005_src0_channel;                                                         // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                           // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                     // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                           // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                   // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [92:0] rsp_xbar_demux_006_src0_data;                                                            // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire  [57:0] rsp_xbar_demux_006_src0_channel;                                                         // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                           // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                     // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                           // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                   // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire  [92:0] rsp_xbar_demux_007_src0_data;                                                            // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire  [57:0] rsp_xbar_demux_007_src0_channel;                                                         // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                           // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                     // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                           // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                   // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	wire  [92:0] rsp_xbar_demux_008_src0_data;                                                            // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	wire  [57:0] rsp_xbar_demux_008_src0_channel;                                                         // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                           // rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                     // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                           // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                   // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	wire  [92:0] rsp_xbar_demux_009_src0_data;                                                            // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	wire  [57:0] rsp_xbar_demux_009_src0_channel;                                                         // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                           // rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                     // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                           // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                   // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux:sink10_startofpacket
	wire  [92:0] rsp_xbar_demux_010_src0_data;                                                            // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux:sink10_data
	wire  [57:0] rsp_xbar_demux_010_src0_channel;                                                         // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                           // rsp_xbar_mux:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                     // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                           // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                   // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux:sink11_startofpacket
	wire  [92:0] rsp_xbar_demux_011_src0_data;                                                            // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux:sink11_data
	wire  [57:0] rsp_xbar_demux_011_src0_channel;                                                         // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                           // rsp_xbar_mux:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                     // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux:sink12_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                           // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux:sink12_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                   // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux:sink12_startofpacket
	wire  [92:0] rsp_xbar_demux_012_src0_data;                                                            // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux:sink12_data
	wire  [57:0] rsp_xbar_demux_012_src0_channel;                                                         // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux:sink12_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                           // rsp_xbar_mux:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                     // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux:sink13_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                           // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux:sink13_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                   // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux:sink13_startofpacket
	wire  [92:0] rsp_xbar_demux_013_src0_data;                                                            // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux:sink13_data
	wire  [57:0] rsp_xbar_demux_013_src0_channel;                                                         // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux:sink13_channel
	wire         rsp_xbar_demux_013_src0_ready;                                                           // rsp_xbar_mux:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire         rsp_xbar_demux_014_src0_endofpacket;                                                     // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux:sink14_endofpacket
	wire         rsp_xbar_demux_014_src0_valid;                                                           // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux:sink14_valid
	wire         rsp_xbar_demux_014_src0_startofpacket;                                                   // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux:sink14_startofpacket
	wire  [92:0] rsp_xbar_demux_014_src0_data;                                                            // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux:sink14_data
	wire  [57:0] rsp_xbar_demux_014_src0_channel;                                                         // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux:sink14_channel
	wire         rsp_xbar_demux_014_src0_ready;                                                           // rsp_xbar_mux:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire         rsp_xbar_demux_015_src0_endofpacket;                                                     // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux:sink15_endofpacket
	wire         rsp_xbar_demux_015_src0_valid;                                                           // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux:sink15_valid
	wire         rsp_xbar_demux_015_src0_startofpacket;                                                   // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux:sink15_startofpacket
	wire  [92:0] rsp_xbar_demux_015_src0_data;                                                            // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux:sink15_data
	wire  [57:0] rsp_xbar_demux_015_src0_channel;                                                         // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux:sink15_channel
	wire         rsp_xbar_demux_015_src0_ready;                                                           // rsp_xbar_mux:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire         rsp_xbar_demux_016_src0_endofpacket;                                                     // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux:sink16_endofpacket
	wire         rsp_xbar_demux_016_src0_valid;                                                           // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux:sink16_valid
	wire         rsp_xbar_demux_016_src0_startofpacket;                                                   // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux:sink16_startofpacket
	wire  [92:0] rsp_xbar_demux_016_src0_data;                                                            // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux:sink16_data
	wire  [57:0] rsp_xbar_demux_016_src0_channel;                                                         // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux:sink16_channel
	wire         rsp_xbar_demux_016_src0_ready;                                                           // rsp_xbar_mux:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire         rsp_xbar_demux_017_src0_endofpacket;                                                     // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux:sink17_endofpacket
	wire         rsp_xbar_demux_017_src0_valid;                                                           // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux:sink17_valid
	wire         rsp_xbar_demux_017_src0_startofpacket;                                                   // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux:sink17_startofpacket
	wire  [92:0] rsp_xbar_demux_017_src0_data;                                                            // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux:sink17_data
	wire  [57:0] rsp_xbar_demux_017_src0_channel;                                                         // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux:sink17_channel
	wire         rsp_xbar_demux_017_src0_ready;                                                           // rsp_xbar_mux:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire         rsp_xbar_demux_018_src0_endofpacket;                                                     // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux:sink18_endofpacket
	wire         rsp_xbar_demux_018_src0_valid;                                                           // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux:sink18_valid
	wire         rsp_xbar_demux_018_src0_startofpacket;                                                   // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux:sink18_startofpacket
	wire  [92:0] rsp_xbar_demux_018_src0_data;                                                            // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux:sink18_data
	wire  [57:0] rsp_xbar_demux_018_src0_channel;                                                         // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux:sink18_channel
	wire         rsp_xbar_demux_018_src0_ready;                                                           // rsp_xbar_mux:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire         rsp_xbar_demux_019_src0_endofpacket;                                                     // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux:sink19_endofpacket
	wire         rsp_xbar_demux_019_src0_valid;                                                           // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux:sink19_valid
	wire         rsp_xbar_demux_019_src0_startofpacket;                                                   // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux:sink19_startofpacket
	wire  [92:0] rsp_xbar_demux_019_src0_data;                                                            // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux:sink19_data
	wire  [57:0] rsp_xbar_demux_019_src0_channel;                                                         // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux:sink19_channel
	wire         rsp_xbar_demux_019_src0_ready;                                                           // rsp_xbar_mux:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire         rsp_xbar_demux_020_src0_endofpacket;                                                     // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux:sink20_endofpacket
	wire         rsp_xbar_demux_020_src0_valid;                                                           // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux:sink20_valid
	wire         rsp_xbar_demux_020_src0_startofpacket;                                                   // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux:sink20_startofpacket
	wire  [92:0] rsp_xbar_demux_020_src0_data;                                                            // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux:sink20_data
	wire  [57:0] rsp_xbar_demux_020_src0_channel;                                                         // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux:sink20_channel
	wire         rsp_xbar_demux_020_src0_ready;                                                           // rsp_xbar_mux:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire         rsp_xbar_demux_021_src0_endofpacket;                                                     // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux:sink21_endofpacket
	wire         rsp_xbar_demux_021_src0_valid;                                                           // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux:sink21_valid
	wire         rsp_xbar_demux_021_src0_startofpacket;                                                   // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux:sink21_startofpacket
	wire  [92:0] rsp_xbar_demux_021_src0_data;                                                            // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux:sink21_data
	wire  [57:0] rsp_xbar_demux_021_src0_channel;                                                         // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux:sink21_channel
	wire         rsp_xbar_demux_021_src0_ready;                                                           // rsp_xbar_mux:sink21_ready -> rsp_xbar_demux_021:src0_ready
	wire         rsp_xbar_demux_022_src0_endofpacket;                                                     // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux:sink22_endofpacket
	wire         rsp_xbar_demux_022_src0_valid;                                                           // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux:sink22_valid
	wire         rsp_xbar_demux_022_src0_startofpacket;                                                   // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux:sink22_startofpacket
	wire  [92:0] rsp_xbar_demux_022_src0_data;                                                            // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux:sink22_data
	wire  [57:0] rsp_xbar_demux_022_src0_channel;                                                         // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux:sink22_channel
	wire         rsp_xbar_demux_022_src0_ready;                                                           // rsp_xbar_mux:sink22_ready -> rsp_xbar_demux_022:src0_ready
	wire         rsp_xbar_demux_023_src0_endofpacket;                                                     // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux:sink23_endofpacket
	wire         rsp_xbar_demux_023_src0_valid;                                                           // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux:sink23_valid
	wire         rsp_xbar_demux_023_src0_startofpacket;                                                   // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux:sink23_startofpacket
	wire  [92:0] rsp_xbar_demux_023_src0_data;                                                            // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux:sink23_data
	wire  [57:0] rsp_xbar_demux_023_src0_channel;                                                         // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux:sink23_channel
	wire         rsp_xbar_demux_023_src0_ready;                                                           // rsp_xbar_mux:sink23_ready -> rsp_xbar_demux_023:src0_ready
	wire         rsp_xbar_demux_024_src0_endofpacket;                                                     // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux:sink24_endofpacket
	wire         rsp_xbar_demux_024_src0_valid;                                                           // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux:sink24_valid
	wire         rsp_xbar_demux_024_src0_startofpacket;                                                   // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux:sink24_startofpacket
	wire  [92:0] rsp_xbar_demux_024_src0_data;                                                            // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux:sink24_data
	wire  [57:0] rsp_xbar_demux_024_src0_channel;                                                         // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux:sink24_channel
	wire         rsp_xbar_demux_024_src0_ready;                                                           // rsp_xbar_mux:sink24_ready -> rsp_xbar_demux_024:src0_ready
	wire         rsp_xbar_demux_025_src0_endofpacket;                                                     // rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux:sink25_endofpacket
	wire         rsp_xbar_demux_025_src0_valid;                                                           // rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux:sink25_valid
	wire         rsp_xbar_demux_025_src0_startofpacket;                                                   // rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux:sink25_startofpacket
	wire  [92:0] rsp_xbar_demux_025_src0_data;                                                            // rsp_xbar_demux_025:src0_data -> rsp_xbar_mux:sink25_data
	wire  [57:0] rsp_xbar_demux_025_src0_channel;                                                         // rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux:sink25_channel
	wire         rsp_xbar_demux_025_src0_ready;                                                           // rsp_xbar_mux:sink25_ready -> rsp_xbar_demux_025:src0_ready
	wire         rsp_xbar_demux_026_src0_endofpacket;                                                     // rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux:sink26_endofpacket
	wire         rsp_xbar_demux_026_src0_valid;                                                           // rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux:sink26_valid
	wire         rsp_xbar_demux_026_src0_startofpacket;                                                   // rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux:sink26_startofpacket
	wire  [92:0] rsp_xbar_demux_026_src0_data;                                                            // rsp_xbar_demux_026:src0_data -> rsp_xbar_mux:sink26_data
	wire  [57:0] rsp_xbar_demux_026_src0_channel;                                                         // rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux:sink26_channel
	wire         rsp_xbar_demux_026_src0_ready;                                                           // rsp_xbar_mux:sink26_ready -> rsp_xbar_demux_026:src0_ready
	wire         rsp_xbar_demux_027_src0_endofpacket;                                                     // rsp_xbar_demux_027:src0_endofpacket -> rsp_xbar_mux:sink27_endofpacket
	wire         rsp_xbar_demux_027_src0_valid;                                                           // rsp_xbar_demux_027:src0_valid -> rsp_xbar_mux:sink27_valid
	wire         rsp_xbar_demux_027_src0_startofpacket;                                                   // rsp_xbar_demux_027:src0_startofpacket -> rsp_xbar_mux:sink27_startofpacket
	wire  [92:0] rsp_xbar_demux_027_src0_data;                                                            // rsp_xbar_demux_027:src0_data -> rsp_xbar_mux:sink27_data
	wire  [57:0] rsp_xbar_demux_027_src0_channel;                                                         // rsp_xbar_demux_027:src0_channel -> rsp_xbar_mux:sink27_channel
	wire         rsp_xbar_demux_027_src0_ready;                                                           // rsp_xbar_mux:sink27_ready -> rsp_xbar_demux_027:src0_ready
	wire         rsp_xbar_demux_028_src0_endofpacket;                                                     // rsp_xbar_demux_028:src0_endofpacket -> rsp_xbar_mux:sink28_endofpacket
	wire         rsp_xbar_demux_028_src0_valid;                                                           // rsp_xbar_demux_028:src0_valid -> rsp_xbar_mux:sink28_valid
	wire         rsp_xbar_demux_028_src0_startofpacket;                                                   // rsp_xbar_demux_028:src0_startofpacket -> rsp_xbar_mux:sink28_startofpacket
	wire  [92:0] rsp_xbar_demux_028_src0_data;                                                            // rsp_xbar_demux_028:src0_data -> rsp_xbar_mux:sink28_data
	wire  [57:0] rsp_xbar_demux_028_src0_channel;                                                         // rsp_xbar_demux_028:src0_channel -> rsp_xbar_mux:sink28_channel
	wire         rsp_xbar_demux_028_src0_ready;                                                           // rsp_xbar_mux:sink28_ready -> rsp_xbar_demux_028:src0_ready
	wire         rsp_xbar_demux_029_src0_endofpacket;                                                     // rsp_xbar_demux_029:src0_endofpacket -> rsp_xbar_mux:sink29_endofpacket
	wire         rsp_xbar_demux_029_src0_valid;                                                           // rsp_xbar_demux_029:src0_valid -> rsp_xbar_mux:sink29_valid
	wire         rsp_xbar_demux_029_src0_startofpacket;                                                   // rsp_xbar_demux_029:src0_startofpacket -> rsp_xbar_mux:sink29_startofpacket
	wire  [92:0] rsp_xbar_demux_029_src0_data;                                                            // rsp_xbar_demux_029:src0_data -> rsp_xbar_mux:sink29_data
	wire  [57:0] rsp_xbar_demux_029_src0_channel;                                                         // rsp_xbar_demux_029:src0_channel -> rsp_xbar_mux:sink29_channel
	wire         rsp_xbar_demux_029_src0_ready;                                                           // rsp_xbar_mux:sink29_ready -> rsp_xbar_demux_029:src0_ready
	wire         rsp_xbar_demux_030_src0_endofpacket;                                                     // rsp_xbar_demux_030:src0_endofpacket -> rsp_xbar_mux:sink30_endofpacket
	wire         rsp_xbar_demux_030_src0_valid;                                                           // rsp_xbar_demux_030:src0_valid -> rsp_xbar_mux:sink30_valid
	wire         rsp_xbar_demux_030_src0_startofpacket;                                                   // rsp_xbar_demux_030:src0_startofpacket -> rsp_xbar_mux:sink30_startofpacket
	wire  [92:0] rsp_xbar_demux_030_src0_data;                                                            // rsp_xbar_demux_030:src0_data -> rsp_xbar_mux:sink30_data
	wire  [57:0] rsp_xbar_demux_030_src0_channel;                                                         // rsp_xbar_demux_030:src0_channel -> rsp_xbar_mux:sink30_channel
	wire         rsp_xbar_demux_030_src0_ready;                                                           // rsp_xbar_mux:sink30_ready -> rsp_xbar_demux_030:src0_ready
	wire         rsp_xbar_demux_031_src0_endofpacket;                                                     // rsp_xbar_demux_031:src0_endofpacket -> rsp_xbar_mux:sink31_endofpacket
	wire         rsp_xbar_demux_031_src0_valid;                                                           // rsp_xbar_demux_031:src0_valid -> rsp_xbar_mux:sink31_valid
	wire         rsp_xbar_demux_031_src0_startofpacket;                                                   // rsp_xbar_demux_031:src0_startofpacket -> rsp_xbar_mux:sink31_startofpacket
	wire  [92:0] rsp_xbar_demux_031_src0_data;                                                            // rsp_xbar_demux_031:src0_data -> rsp_xbar_mux:sink31_data
	wire  [57:0] rsp_xbar_demux_031_src0_channel;                                                         // rsp_xbar_demux_031:src0_channel -> rsp_xbar_mux:sink31_channel
	wire         rsp_xbar_demux_031_src0_ready;                                                           // rsp_xbar_mux:sink31_ready -> rsp_xbar_demux_031:src0_ready
	wire         rsp_xbar_demux_032_src0_endofpacket;                                                     // rsp_xbar_demux_032:src0_endofpacket -> rsp_xbar_mux:sink32_endofpacket
	wire         rsp_xbar_demux_032_src0_valid;                                                           // rsp_xbar_demux_032:src0_valid -> rsp_xbar_mux:sink32_valid
	wire         rsp_xbar_demux_032_src0_startofpacket;                                                   // rsp_xbar_demux_032:src0_startofpacket -> rsp_xbar_mux:sink32_startofpacket
	wire  [92:0] rsp_xbar_demux_032_src0_data;                                                            // rsp_xbar_demux_032:src0_data -> rsp_xbar_mux:sink32_data
	wire  [57:0] rsp_xbar_demux_032_src0_channel;                                                         // rsp_xbar_demux_032:src0_channel -> rsp_xbar_mux:sink32_channel
	wire         rsp_xbar_demux_032_src0_ready;                                                           // rsp_xbar_mux:sink32_ready -> rsp_xbar_demux_032:src0_ready
	wire         rsp_xbar_demux_033_src0_endofpacket;                                                     // rsp_xbar_demux_033:src0_endofpacket -> rsp_xbar_mux:sink33_endofpacket
	wire         rsp_xbar_demux_033_src0_valid;                                                           // rsp_xbar_demux_033:src0_valid -> rsp_xbar_mux:sink33_valid
	wire         rsp_xbar_demux_033_src0_startofpacket;                                                   // rsp_xbar_demux_033:src0_startofpacket -> rsp_xbar_mux:sink33_startofpacket
	wire  [92:0] rsp_xbar_demux_033_src0_data;                                                            // rsp_xbar_demux_033:src0_data -> rsp_xbar_mux:sink33_data
	wire  [57:0] rsp_xbar_demux_033_src0_channel;                                                         // rsp_xbar_demux_033:src0_channel -> rsp_xbar_mux:sink33_channel
	wire         rsp_xbar_demux_033_src0_ready;                                                           // rsp_xbar_mux:sink33_ready -> rsp_xbar_demux_033:src0_ready
	wire         rsp_xbar_demux_034_src0_endofpacket;                                                     // rsp_xbar_demux_034:src0_endofpacket -> rsp_xbar_mux:sink34_endofpacket
	wire         rsp_xbar_demux_034_src0_valid;                                                           // rsp_xbar_demux_034:src0_valid -> rsp_xbar_mux:sink34_valid
	wire         rsp_xbar_demux_034_src0_startofpacket;                                                   // rsp_xbar_demux_034:src0_startofpacket -> rsp_xbar_mux:sink34_startofpacket
	wire  [92:0] rsp_xbar_demux_034_src0_data;                                                            // rsp_xbar_demux_034:src0_data -> rsp_xbar_mux:sink34_data
	wire  [57:0] rsp_xbar_demux_034_src0_channel;                                                         // rsp_xbar_demux_034:src0_channel -> rsp_xbar_mux:sink34_channel
	wire         rsp_xbar_demux_034_src0_ready;                                                           // rsp_xbar_mux:sink34_ready -> rsp_xbar_demux_034:src0_ready
	wire         rsp_xbar_demux_035_src0_endofpacket;                                                     // rsp_xbar_demux_035:src0_endofpacket -> rsp_xbar_mux:sink35_endofpacket
	wire         rsp_xbar_demux_035_src0_valid;                                                           // rsp_xbar_demux_035:src0_valid -> rsp_xbar_mux:sink35_valid
	wire         rsp_xbar_demux_035_src0_startofpacket;                                                   // rsp_xbar_demux_035:src0_startofpacket -> rsp_xbar_mux:sink35_startofpacket
	wire  [92:0] rsp_xbar_demux_035_src0_data;                                                            // rsp_xbar_demux_035:src0_data -> rsp_xbar_mux:sink35_data
	wire  [57:0] rsp_xbar_demux_035_src0_channel;                                                         // rsp_xbar_demux_035:src0_channel -> rsp_xbar_mux:sink35_channel
	wire         rsp_xbar_demux_035_src0_ready;                                                           // rsp_xbar_mux:sink35_ready -> rsp_xbar_demux_035:src0_ready
	wire         rsp_xbar_demux_036_src0_endofpacket;                                                     // rsp_xbar_demux_036:src0_endofpacket -> rsp_xbar_mux:sink36_endofpacket
	wire         rsp_xbar_demux_036_src0_valid;                                                           // rsp_xbar_demux_036:src0_valid -> rsp_xbar_mux:sink36_valid
	wire         rsp_xbar_demux_036_src0_startofpacket;                                                   // rsp_xbar_demux_036:src0_startofpacket -> rsp_xbar_mux:sink36_startofpacket
	wire  [92:0] rsp_xbar_demux_036_src0_data;                                                            // rsp_xbar_demux_036:src0_data -> rsp_xbar_mux:sink36_data
	wire  [57:0] rsp_xbar_demux_036_src0_channel;                                                         // rsp_xbar_demux_036:src0_channel -> rsp_xbar_mux:sink36_channel
	wire         rsp_xbar_demux_036_src0_ready;                                                           // rsp_xbar_mux:sink36_ready -> rsp_xbar_demux_036:src0_ready
	wire         rsp_xbar_demux_037_src0_endofpacket;                                                     // rsp_xbar_demux_037:src0_endofpacket -> rsp_xbar_mux:sink37_endofpacket
	wire         rsp_xbar_demux_037_src0_valid;                                                           // rsp_xbar_demux_037:src0_valid -> rsp_xbar_mux:sink37_valid
	wire         rsp_xbar_demux_037_src0_startofpacket;                                                   // rsp_xbar_demux_037:src0_startofpacket -> rsp_xbar_mux:sink37_startofpacket
	wire  [92:0] rsp_xbar_demux_037_src0_data;                                                            // rsp_xbar_demux_037:src0_data -> rsp_xbar_mux:sink37_data
	wire  [57:0] rsp_xbar_demux_037_src0_channel;                                                         // rsp_xbar_demux_037:src0_channel -> rsp_xbar_mux:sink37_channel
	wire         rsp_xbar_demux_037_src0_ready;                                                           // rsp_xbar_mux:sink37_ready -> rsp_xbar_demux_037:src0_ready
	wire         rsp_xbar_demux_038_src0_endofpacket;                                                     // rsp_xbar_demux_038:src0_endofpacket -> rsp_xbar_mux:sink38_endofpacket
	wire         rsp_xbar_demux_038_src0_valid;                                                           // rsp_xbar_demux_038:src0_valid -> rsp_xbar_mux:sink38_valid
	wire         rsp_xbar_demux_038_src0_startofpacket;                                                   // rsp_xbar_demux_038:src0_startofpacket -> rsp_xbar_mux:sink38_startofpacket
	wire  [92:0] rsp_xbar_demux_038_src0_data;                                                            // rsp_xbar_demux_038:src0_data -> rsp_xbar_mux:sink38_data
	wire  [57:0] rsp_xbar_demux_038_src0_channel;                                                         // rsp_xbar_demux_038:src0_channel -> rsp_xbar_mux:sink38_channel
	wire         rsp_xbar_demux_038_src0_ready;                                                           // rsp_xbar_mux:sink38_ready -> rsp_xbar_demux_038:src0_ready
	wire         rsp_xbar_demux_039_src0_endofpacket;                                                     // rsp_xbar_demux_039:src0_endofpacket -> rsp_xbar_mux:sink39_endofpacket
	wire         rsp_xbar_demux_039_src0_valid;                                                           // rsp_xbar_demux_039:src0_valid -> rsp_xbar_mux:sink39_valid
	wire         rsp_xbar_demux_039_src0_startofpacket;                                                   // rsp_xbar_demux_039:src0_startofpacket -> rsp_xbar_mux:sink39_startofpacket
	wire  [92:0] rsp_xbar_demux_039_src0_data;                                                            // rsp_xbar_demux_039:src0_data -> rsp_xbar_mux:sink39_data
	wire  [57:0] rsp_xbar_demux_039_src0_channel;                                                         // rsp_xbar_demux_039:src0_channel -> rsp_xbar_mux:sink39_channel
	wire         rsp_xbar_demux_039_src0_ready;                                                           // rsp_xbar_mux:sink39_ready -> rsp_xbar_demux_039:src0_ready
	wire         rsp_xbar_demux_040_src0_endofpacket;                                                     // rsp_xbar_demux_040:src0_endofpacket -> rsp_xbar_mux:sink40_endofpacket
	wire         rsp_xbar_demux_040_src0_valid;                                                           // rsp_xbar_demux_040:src0_valid -> rsp_xbar_mux:sink40_valid
	wire         rsp_xbar_demux_040_src0_startofpacket;                                                   // rsp_xbar_demux_040:src0_startofpacket -> rsp_xbar_mux:sink40_startofpacket
	wire  [92:0] rsp_xbar_demux_040_src0_data;                                                            // rsp_xbar_demux_040:src0_data -> rsp_xbar_mux:sink40_data
	wire  [57:0] rsp_xbar_demux_040_src0_channel;                                                         // rsp_xbar_demux_040:src0_channel -> rsp_xbar_mux:sink40_channel
	wire         rsp_xbar_demux_040_src0_ready;                                                           // rsp_xbar_mux:sink40_ready -> rsp_xbar_demux_040:src0_ready
	wire         rsp_xbar_demux_041_src0_endofpacket;                                                     // rsp_xbar_demux_041:src0_endofpacket -> rsp_xbar_mux:sink41_endofpacket
	wire         rsp_xbar_demux_041_src0_valid;                                                           // rsp_xbar_demux_041:src0_valid -> rsp_xbar_mux:sink41_valid
	wire         rsp_xbar_demux_041_src0_startofpacket;                                                   // rsp_xbar_demux_041:src0_startofpacket -> rsp_xbar_mux:sink41_startofpacket
	wire  [92:0] rsp_xbar_demux_041_src0_data;                                                            // rsp_xbar_demux_041:src0_data -> rsp_xbar_mux:sink41_data
	wire  [57:0] rsp_xbar_demux_041_src0_channel;                                                         // rsp_xbar_demux_041:src0_channel -> rsp_xbar_mux:sink41_channel
	wire         rsp_xbar_demux_041_src0_ready;                                                           // rsp_xbar_mux:sink41_ready -> rsp_xbar_demux_041:src0_ready
	wire         rsp_xbar_demux_042_src0_endofpacket;                                                     // rsp_xbar_demux_042:src0_endofpacket -> rsp_xbar_mux:sink42_endofpacket
	wire         rsp_xbar_demux_042_src0_valid;                                                           // rsp_xbar_demux_042:src0_valid -> rsp_xbar_mux:sink42_valid
	wire         rsp_xbar_demux_042_src0_startofpacket;                                                   // rsp_xbar_demux_042:src0_startofpacket -> rsp_xbar_mux:sink42_startofpacket
	wire  [92:0] rsp_xbar_demux_042_src0_data;                                                            // rsp_xbar_demux_042:src0_data -> rsp_xbar_mux:sink42_data
	wire  [57:0] rsp_xbar_demux_042_src0_channel;                                                         // rsp_xbar_demux_042:src0_channel -> rsp_xbar_mux:sink42_channel
	wire         rsp_xbar_demux_042_src0_ready;                                                           // rsp_xbar_mux:sink42_ready -> rsp_xbar_demux_042:src0_ready
	wire         rsp_xbar_demux_043_src0_endofpacket;                                                     // rsp_xbar_demux_043:src0_endofpacket -> rsp_xbar_mux:sink43_endofpacket
	wire         rsp_xbar_demux_043_src0_valid;                                                           // rsp_xbar_demux_043:src0_valid -> rsp_xbar_mux:sink43_valid
	wire         rsp_xbar_demux_043_src0_startofpacket;                                                   // rsp_xbar_demux_043:src0_startofpacket -> rsp_xbar_mux:sink43_startofpacket
	wire  [92:0] rsp_xbar_demux_043_src0_data;                                                            // rsp_xbar_demux_043:src0_data -> rsp_xbar_mux:sink43_data
	wire  [57:0] rsp_xbar_demux_043_src0_channel;                                                         // rsp_xbar_demux_043:src0_channel -> rsp_xbar_mux:sink43_channel
	wire         rsp_xbar_demux_043_src0_ready;                                                           // rsp_xbar_mux:sink43_ready -> rsp_xbar_demux_043:src0_ready
	wire         rsp_xbar_demux_044_src0_endofpacket;                                                     // rsp_xbar_demux_044:src0_endofpacket -> rsp_xbar_mux:sink44_endofpacket
	wire         rsp_xbar_demux_044_src0_valid;                                                           // rsp_xbar_demux_044:src0_valid -> rsp_xbar_mux:sink44_valid
	wire         rsp_xbar_demux_044_src0_startofpacket;                                                   // rsp_xbar_demux_044:src0_startofpacket -> rsp_xbar_mux:sink44_startofpacket
	wire  [92:0] rsp_xbar_demux_044_src0_data;                                                            // rsp_xbar_demux_044:src0_data -> rsp_xbar_mux:sink44_data
	wire  [57:0] rsp_xbar_demux_044_src0_channel;                                                         // rsp_xbar_demux_044:src0_channel -> rsp_xbar_mux:sink44_channel
	wire         rsp_xbar_demux_044_src0_ready;                                                           // rsp_xbar_mux:sink44_ready -> rsp_xbar_demux_044:src0_ready
	wire         rsp_xbar_demux_045_src0_endofpacket;                                                     // rsp_xbar_demux_045:src0_endofpacket -> rsp_xbar_mux:sink45_endofpacket
	wire         rsp_xbar_demux_045_src0_valid;                                                           // rsp_xbar_demux_045:src0_valid -> rsp_xbar_mux:sink45_valid
	wire         rsp_xbar_demux_045_src0_startofpacket;                                                   // rsp_xbar_demux_045:src0_startofpacket -> rsp_xbar_mux:sink45_startofpacket
	wire  [92:0] rsp_xbar_demux_045_src0_data;                                                            // rsp_xbar_demux_045:src0_data -> rsp_xbar_mux:sink45_data
	wire  [57:0] rsp_xbar_demux_045_src0_channel;                                                         // rsp_xbar_demux_045:src0_channel -> rsp_xbar_mux:sink45_channel
	wire         rsp_xbar_demux_045_src0_ready;                                                           // rsp_xbar_mux:sink45_ready -> rsp_xbar_demux_045:src0_ready
	wire         rsp_xbar_demux_046_src0_endofpacket;                                                     // rsp_xbar_demux_046:src0_endofpacket -> rsp_xbar_mux:sink46_endofpacket
	wire         rsp_xbar_demux_046_src0_valid;                                                           // rsp_xbar_demux_046:src0_valid -> rsp_xbar_mux:sink46_valid
	wire         rsp_xbar_demux_046_src0_startofpacket;                                                   // rsp_xbar_demux_046:src0_startofpacket -> rsp_xbar_mux:sink46_startofpacket
	wire  [92:0] rsp_xbar_demux_046_src0_data;                                                            // rsp_xbar_demux_046:src0_data -> rsp_xbar_mux:sink46_data
	wire  [57:0] rsp_xbar_demux_046_src0_channel;                                                         // rsp_xbar_demux_046:src0_channel -> rsp_xbar_mux:sink46_channel
	wire         rsp_xbar_demux_046_src0_ready;                                                           // rsp_xbar_mux:sink46_ready -> rsp_xbar_demux_046:src0_ready
	wire         rsp_xbar_demux_047_src0_endofpacket;                                                     // rsp_xbar_demux_047:src0_endofpacket -> rsp_xbar_mux:sink47_endofpacket
	wire         rsp_xbar_demux_047_src0_valid;                                                           // rsp_xbar_demux_047:src0_valid -> rsp_xbar_mux:sink47_valid
	wire         rsp_xbar_demux_047_src0_startofpacket;                                                   // rsp_xbar_demux_047:src0_startofpacket -> rsp_xbar_mux:sink47_startofpacket
	wire  [92:0] rsp_xbar_demux_047_src0_data;                                                            // rsp_xbar_demux_047:src0_data -> rsp_xbar_mux:sink47_data
	wire  [57:0] rsp_xbar_demux_047_src0_channel;                                                         // rsp_xbar_demux_047:src0_channel -> rsp_xbar_mux:sink47_channel
	wire         rsp_xbar_demux_047_src0_ready;                                                           // rsp_xbar_mux:sink47_ready -> rsp_xbar_demux_047:src0_ready
	wire         rsp_xbar_demux_048_src0_endofpacket;                                                     // rsp_xbar_demux_048:src0_endofpacket -> rsp_xbar_mux:sink48_endofpacket
	wire         rsp_xbar_demux_048_src0_valid;                                                           // rsp_xbar_demux_048:src0_valid -> rsp_xbar_mux:sink48_valid
	wire         rsp_xbar_demux_048_src0_startofpacket;                                                   // rsp_xbar_demux_048:src0_startofpacket -> rsp_xbar_mux:sink48_startofpacket
	wire  [92:0] rsp_xbar_demux_048_src0_data;                                                            // rsp_xbar_demux_048:src0_data -> rsp_xbar_mux:sink48_data
	wire  [57:0] rsp_xbar_demux_048_src0_channel;                                                         // rsp_xbar_demux_048:src0_channel -> rsp_xbar_mux:sink48_channel
	wire         rsp_xbar_demux_048_src0_ready;                                                           // rsp_xbar_mux:sink48_ready -> rsp_xbar_demux_048:src0_ready
	wire         rsp_xbar_demux_049_src0_endofpacket;                                                     // rsp_xbar_demux_049:src0_endofpacket -> rsp_xbar_mux:sink49_endofpacket
	wire         rsp_xbar_demux_049_src0_valid;                                                           // rsp_xbar_demux_049:src0_valid -> rsp_xbar_mux:sink49_valid
	wire         rsp_xbar_demux_049_src0_startofpacket;                                                   // rsp_xbar_demux_049:src0_startofpacket -> rsp_xbar_mux:sink49_startofpacket
	wire  [92:0] rsp_xbar_demux_049_src0_data;                                                            // rsp_xbar_demux_049:src0_data -> rsp_xbar_mux:sink49_data
	wire  [57:0] rsp_xbar_demux_049_src0_channel;                                                         // rsp_xbar_demux_049:src0_channel -> rsp_xbar_mux:sink49_channel
	wire         rsp_xbar_demux_049_src0_ready;                                                           // rsp_xbar_mux:sink49_ready -> rsp_xbar_demux_049:src0_ready
	wire         rsp_xbar_demux_050_src0_endofpacket;                                                     // rsp_xbar_demux_050:src0_endofpacket -> rsp_xbar_mux:sink50_endofpacket
	wire         rsp_xbar_demux_050_src0_valid;                                                           // rsp_xbar_demux_050:src0_valid -> rsp_xbar_mux:sink50_valid
	wire         rsp_xbar_demux_050_src0_startofpacket;                                                   // rsp_xbar_demux_050:src0_startofpacket -> rsp_xbar_mux:sink50_startofpacket
	wire  [92:0] rsp_xbar_demux_050_src0_data;                                                            // rsp_xbar_demux_050:src0_data -> rsp_xbar_mux:sink50_data
	wire  [57:0] rsp_xbar_demux_050_src0_channel;                                                         // rsp_xbar_demux_050:src0_channel -> rsp_xbar_mux:sink50_channel
	wire         rsp_xbar_demux_050_src0_ready;                                                           // rsp_xbar_mux:sink50_ready -> rsp_xbar_demux_050:src0_ready
	wire         rsp_xbar_demux_051_src0_endofpacket;                                                     // rsp_xbar_demux_051:src0_endofpacket -> rsp_xbar_mux:sink51_endofpacket
	wire         rsp_xbar_demux_051_src0_valid;                                                           // rsp_xbar_demux_051:src0_valid -> rsp_xbar_mux:sink51_valid
	wire         rsp_xbar_demux_051_src0_startofpacket;                                                   // rsp_xbar_demux_051:src0_startofpacket -> rsp_xbar_mux:sink51_startofpacket
	wire  [92:0] rsp_xbar_demux_051_src0_data;                                                            // rsp_xbar_demux_051:src0_data -> rsp_xbar_mux:sink51_data
	wire  [57:0] rsp_xbar_demux_051_src0_channel;                                                         // rsp_xbar_demux_051:src0_channel -> rsp_xbar_mux:sink51_channel
	wire         rsp_xbar_demux_051_src0_ready;                                                           // rsp_xbar_mux:sink51_ready -> rsp_xbar_demux_051:src0_ready
	wire         rsp_xbar_demux_052_src0_endofpacket;                                                     // rsp_xbar_demux_052:src0_endofpacket -> rsp_xbar_mux:sink52_endofpacket
	wire         rsp_xbar_demux_052_src0_valid;                                                           // rsp_xbar_demux_052:src0_valid -> rsp_xbar_mux:sink52_valid
	wire         rsp_xbar_demux_052_src0_startofpacket;                                                   // rsp_xbar_demux_052:src0_startofpacket -> rsp_xbar_mux:sink52_startofpacket
	wire  [92:0] rsp_xbar_demux_052_src0_data;                                                            // rsp_xbar_demux_052:src0_data -> rsp_xbar_mux:sink52_data
	wire  [57:0] rsp_xbar_demux_052_src0_channel;                                                         // rsp_xbar_demux_052:src0_channel -> rsp_xbar_mux:sink52_channel
	wire         rsp_xbar_demux_052_src0_ready;                                                           // rsp_xbar_mux:sink52_ready -> rsp_xbar_demux_052:src0_ready
	wire         rsp_xbar_demux_053_src0_endofpacket;                                                     // rsp_xbar_demux_053:src0_endofpacket -> rsp_xbar_mux:sink53_endofpacket
	wire         rsp_xbar_demux_053_src0_valid;                                                           // rsp_xbar_demux_053:src0_valid -> rsp_xbar_mux:sink53_valid
	wire         rsp_xbar_demux_053_src0_startofpacket;                                                   // rsp_xbar_demux_053:src0_startofpacket -> rsp_xbar_mux:sink53_startofpacket
	wire  [92:0] rsp_xbar_demux_053_src0_data;                                                            // rsp_xbar_demux_053:src0_data -> rsp_xbar_mux:sink53_data
	wire  [57:0] rsp_xbar_demux_053_src0_channel;                                                         // rsp_xbar_demux_053:src0_channel -> rsp_xbar_mux:sink53_channel
	wire         rsp_xbar_demux_053_src0_ready;                                                           // rsp_xbar_mux:sink53_ready -> rsp_xbar_demux_053:src0_ready
	wire         rsp_xbar_demux_054_src0_endofpacket;                                                     // rsp_xbar_demux_054:src0_endofpacket -> rsp_xbar_mux:sink54_endofpacket
	wire         rsp_xbar_demux_054_src0_valid;                                                           // rsp_xbar_demux_054:src0_valid -> rsp_xbar_mux:sink54_valid
	wire         rsp_xbar_demux_054_src0_startofpacket;                                                   // rsp_xbar_demux_054:src0_startofpacket -> rsp_xbar_mux:sink54_startofpacket
	wire  [92:0] rsp_xbar_demux_054_src0_data;                                                            // rsp_xbar_demux_054:src0_data -> rsp_xbar_mux:sink54_data
	wire  [57:0] rsp_xbar_demux_054_src0_channel;                                                         // rsp_xbar_demux_054:src0_channel -> rsp_xbar_mux:sink54_channel
	wire         rsp_xbar_demux_054_src0_ready;                                                           // rsp_xbar_mux:sink54_ready -> rsp_xbar_demux_054:src0_ready
	wire         rsp_xbar_demux_055_src0_endofpacket;                                                     // rsp_xbar_demux_055:src0_endofpacket -> rsp_xbar_mux:sink55_endofpacket
	wire         rsp_xbar_demux_055_src0_valid;                                                           // rsp_xbar_demux_055:src0_valid -> rsp_xbar_mux:sink55_valid
	wire         rsp_xbar_demux_055_src0_startofpacket;                                                   // rsp_xbar_demux_055:src0_startofpacket -> rsp_xbar_mux:sink55_startofpacket
	wire  [92:0] rsp_xbar_demux_055_src0_data;                                                            // rsp_xbar_demux_055:src0_data -> rsp_xbar_mux:sink55_data
	wire  [57:0] rsp_xbar_demux_055_src0_channel;                                                         // rsp_xbar_demux_055:src0_channel -> rsp_xbar_mux:sink55_channel
	wire         rsp_xbar_demux_055_src0_ready;                                                           // rsp_xbar_mux:sink55_ready -> rsp_xbar_demux_055:src0_ready
	wire         rsp_xbar_demux_056_src0_endofpacket;                                                     // rsp_xbar_demux_056:src0_endofpacket -> rsp_xbar_mux:sink56_endofpacket
	wire         rsp_xbar_demux_056_src0_valid;                                                           // rsp_xbar_demux_056:src0_valid -> rsp_xbar_mux:sink56_valid
	wire         rsp_xbar_demux_056_src0_startofpacket;                                                   // rsp_xbar_demux_056:src0_startofpacket -> rsp_xbar_mux:sink56_startofpacket
	wire  [92:0] rsp_xbar_demux_056_src0_data;                                                            // rsp_xbar_demux_056:src0_data -> rsp_xbar_mux:sink56_data
	wire  [57:0] rsp_xbar_demux_056_src0_channel;                                                         // rsp_xbar_demux_056:src0_channel -> rsp_xbar_mux:sink56_channel
	wire         rsp_xbar_demux_056_src0_ready;                                                           // rsp_xbar_mux:sink56_ready -> rsp_xbar_demux_056:src0_ready
	wire         rsp_xbar_demux_057_src0_endofpacket;                                                     // rsp_xbar_demux_057:src0_endofpacket -> rsp_xbar_mux:sink57_endofpacket
	wire         rsp_xbar_demux_057_src0_valid;                                                           // rsp_xbar_demux_057:src0_valid -> rsp_xbar_mux:sink57_valid
	wire         rsp_xbar_demux_057_src0_startofpacket;                                                   // rsp_xbar_demux_057:src0_startofpacket -> rsp_xbar_mux:sink57_startofpacket
	wire  [92:0] rsp_xbar_demux_057_src0_data;                                                            // rsp_xbar_demux_057:src0_data -> rsp_xbar_mux:sink57_data
	wire  [57:0] rsp_xbar_demux_057_src0_channel;                                                         // rsp_xbar_demux_057:src0_channel -> rsp_xbar_mux:sink57_channel
	wire         rsp_xbar_demux_057_src0_ready;                                                           // rsp_xbar_mux:sink57_ready -> rsp_xbar_demux_057:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                             // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                           // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [92:0] limiter_cmd_src_data;                                                                    // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire  [57:0] limiter_cmd_src_channel;                                                                 // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                   // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                            // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                  // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                          // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [92:0] rsp_xbar_mux_src_data;                                                                   // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire  [57:0] rsp_xbar_mux_src_channel;                                                                // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                  // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         cmd_xbar_demux_src0_ready;                                                               // SysID_SysID_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire         id_router_src_endofpacket;                                                               // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                     // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                             // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [92:0] id_router_src_data;                                                                      // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [57:0] id_router_src_channel;                                                                   // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                     // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_demux_src1_ready;                                                               // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire         id_router_001_src_endofpacket;                                                           // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                 // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                         // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [92:0] id_router_001_src_data;                                                                  // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [57:0] id_router_001_src_channel;                                                               // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                 // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_src2_ready;                                                               // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	wire         id_router_002_src_endofpacket;                                                           // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                 // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                         // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [92:0] id_router_002_src_data;                                                                  // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [57:0] id_router_002_src_channel;                                                               // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                 // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_src3_ready;                                                               // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src3_ready
	wire         id_router_003_src_endofpacket;                                                           // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                 // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                         // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [92:0] id_router_003_src_data;                                                                  // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [57:0] id_router_003_src_channel;                                                               // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                 // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_src4_ready;                                                               // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src4_ready
	wire         id_router_004_src_endofpacket;                                                           // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                 // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                         // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [92:0] id_router_004_src_data;                                                                  // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [57:0] id_router_004_src_channel;                                                               // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                 // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_src5_ready;                                                               // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src5_ready
	wire         id_router_005_src_endofpacket;                                                           // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                 // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                         // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [92:0] id_router_005_src_data;                                                                  // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [57:0] id_router_005_src_channel;                                                               // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                 // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_src6_ready;                                                               // width_adapter:in_ready -> cmd_xbar_demux:src6_ready
	wire         width_adapter_src_endofpacket;                                                           // width_adapter:out_endofpacket -> burst_adapter_005:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                 // width_adapter:out_valid -> burst_adapter_005:sink0_valid
	wire         width_adapter_src_startofpacket;                                                         // width_adapter:out_startofpacket -> burst_adapter_005:sink0_startofpacket
	wire  [65:0] width_adapter_src_data;                                                                  // width_adapter:out_data -> burst_adapter_005:sink0_data
	wire         width_adapter_src_ready;                                                                 // burst_adapter_005:sink0_ready -> width_adapter:out_ready
	wire  [57:0] width_adapter_src_channel;                                                               // width_adapter:out_channel -> burst_adapter_005:sink0_channel
	wire         id_router_006_src_endofpacket;                                                           // id_router_006:src_endofpacket -> width_adapter_001:in_endofpacket
	wire         id_router_006_src_valid;                                                                 // id_router_006:src_valid -> width_adapter_001:in_valid
	wire         id_router_006_src_startofpacket;                                                         // id_router_006:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [65:0] id_router_006_src_data;                                                                  // id_router_006:src_data -> width_adapter_001:in_data
	wire  [57:0] id_router_006_src_channel;                                                               // id_router_006:src_channel -> width_adapter_001:in_channel
	wire         id_router_006_src_ready;                                                                 // width_adapter_001:in_ready -> id_router_006:src_ready
	wire         width_adapter_001_src_endofpacket;                                                       // width_adapter_001:out_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         width_adapter_001_src_valid;                                                             // width_adapter_001:out_valid -> rsp_xbar_demux_006:sink_valid
	wire         width_adapter_001_src_startofpacket;                                                     // width_adapter_001:out_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [92:0] width_adapter_001_src_data;                                                              // width_adapter_001:out_data -> rsp_xbar_demux_006:sink_data
	wire         width_adapter_001_src_ready;                                                             // rsp_xbar_demux_006:sink_ready -> width_adapter_001:out_ready
	wire  [57:0] width_adapter_001_src_channel;                                                           // width_adapter_001:out_channel -> rsp_xbar_demux_006:sink_channel
	wire         cmd_xbar_demux_src7_ready;                                                               // width_adapter_002:in_ready -> cmd_xbar_demux:src7_ready
	wire         width_adapter_002_src_endofpacket;                                                       // width_adapter_002:out_endofpacket -> burst_adapter_004:sink0_endofpacket
	wire         width_adapter_002_src_valid;                                                             // width_adapter_002:out_valid -> burst_adapter_004:sink0_valid
	wire         width_adapter_002_src_startofpacket;                                                     // width_adapter_002:out_startofpacket -> burst_adapter_004:sink0_startofpacket
	wire  [65:0] width_adapter_002_src_data;                                                              // width_adapter_002:out_data -> burst_adapter_004:sink0_data
	wire         width_adapter_002_src_ready;                                                             // burst_adapter_004:sink0_ready -> width_adapter_002:out_ready
	wire  [57:0] width_adapter_002_src_channel;                                                           // width_adapter_002:out_channel -> burst_adapter_004:sink0_channel
	wire         id_router_007_src_endofpacket;                                                           // id_router_007:src_endofpacket -> width_adapter_003:in_endofpacket
	wire         id_router_007_src_valid;                                                                 // id_router_007:src_valid -> width_adapter_003:in_valid
	wire         id_router_007_src_startofpacket;                                                         // id_router_007:src_startofpacket -> width_adapter_003:in_startofpacket
	wire  [65:0] id_router_007_src_data;                                                                  // id_router_007:src_data -> width_adapter_003:in_data
	wire  [57:0] id_router_007_src_channel;                                                               // id_router_007:src_channel -> width_adapter_003:in_channel
	wire         id_router_007_src_ready;                                                                 // width_adapter_003:in_ready -> id_router_007:src_ready
	wire         width_adapter_003_src_endofpacket;                                                       // width_adapter_003:out_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         width_adapter_003_src_valid;                                                             // width_adapter_003:out_valid -> rsp_xbar_demux_007:sink_valid
	wire         width_adapter_003_src_startofpacket;                                                     // width_adapter_003:out_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [92:0] width_adapter_003_src_data;                                                              // width_adapter_003:out_data -> rsp_xbar_demux_007:sink_data
	wire         width_adapter_003_src_ready;                                                             // rsp_xbar_demux_007:sink_ready -> width_adapter_003:out_ready
	wire  [57:0] width_adapter_003_src_channel;                                                           // width_adapter_003:out_channel -> rsp_xbar_demux_007:sink_channel
	wire         cmd_xbar_demux_src8_ready;                                                               // width_adapter_004:in_ready -> cmd_xbar_demux:src8_ready
	wire         width_adapter_004_src_endofpacket;                                                       // width_adapter_004:out_endofpacket -> burst_adapter_048:sink0_endofpacket
	wire         width_adapter_004_src_valid;                                                             // width_adapter_004:out_valid -> burst_adapter_048:sink0_valid
	wire         width_adapter_004_src_startofpacket;                                                     // width_adapter_004:out_startofpacket -> burst_adapter_048:sink0_startofpacket
	wire  [65:0] width_adapter_004_src_data;                                                              // width_adapter_004:out_data -> burst_adapter_048:sink0_data
	wire         width_adapter_004_src_ready;                                                             // burst_adapter_048:sink0_ready -> width_adapter_004:out_ready
	wire  [57:0] width_adapter_004_src_channel;                                                           // width_adapter_004:out_channel -> burst_adapter_048:sink0_channel
	wire         id_router_008_src_endofpacket;                                                           // id_router_008:src_endofpacket -> width_adapter_005:in_endofpacket
	wire         id_router_008_src_valid;                                                                 // id_router_008:src_valid -> width_adapter_005:in_valid
	wire         id_router_008_src_startofpacket;                                                         // id_router_008:src_startofpacket -> width_adapter_005:in_startofpacket
	wire  [65:0] id_router_008_src_data;                                                                  // id_router_008:src_data -> width_adapter_005:in_data
	wire  [57:0] id_router_008_src_channel;                                                               // id_router_008:src_channel -> width_adapter_005:in_channel
	wire         id_router_008_src_ready;                                                                 // width_adapter_005:in_ready -> id_router_008:src_ready
	wire         width_adapter_005_src_endofpacket;                                                       // width_adapter_005:out_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         width_adapter_005_src_valid;                                                             // width_adapter_005:out_valid -> rsp_xbar_demux_008:sink_valid
	wire         width_adapter_005_src_startofpacket;                                                     // width_adapter_005:out_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [92:0] width_adapter_005_src_data;                                                              // width_adapter_005:out_data -> rsp_xbar_demux_008:sink_data
	wire         width_adapter_005_src_ready;                                                             // rsp_xbar_demux_008:sink_ready -> width_adapter_005:out_ready
	wire  [57:0] width_adapter_005_src_channel;                                                           // width_adapter_005:out_channel -> rsp_xbar_demux_008:sink_channel
	wire         cmd_xbar_demux_src9_ready;                                                               // width_adapter_006:in_ready -> cmd_xbar_demux:src9_ready
	wire         width_adapter_006_src_endofpacket;                                                       // width_adapter_006:out_endofpacket -> burst_adapter_025:sink0_endofpacket
	wire         width_adapter_006_src_valid;                                                             // width_adapter_006:out_valid -> burst_adapter_025:sink0_valid
	wire         width_adapter_006_src_startofpacket;                                                     // width_adapter_006:out_startofpacket -> burst_adapter_025:sink0_startofpacket
	wire  [65:0] width_adapter_006_src_data;                                                              // width_adapter_006:out_data -> burst_adapter_025:sink0_data
	wire         width_adapter_006_src_ready;                                                             // burst_adapter_025:sink0_ready -> width_adapter_006:out_ready
	wire  [57:0] width_adapter_006_src_channel;                                                           // width_adapter_006:out_channel -> burst_adapter_025:sink0_channel
	wire         id_router_009_src_endofpacket;                                                           // id_router_009:src_endofpacket -> width_adapter_007:in_endofpacket
	wire         id_router_009_src_valid;                                                                 // id_router_009:src_valid -> width_adapter_007:in_valid
	wire         id_router_009_src_startofpacket;                                                         // id_router_009:src_startofpacket -> width_adapter_007:in_startofpacket
	wire  [65:0] id_router_009_src_data;                                                                  // id_router_009:src_data -> width_adapter_007:in_data
	wire  [57:0] id_router_009_src_channel;                                                               // id_router_009:src_channel -> width_adapter_007:in_channel
	wire         id_router_009_src_ready;                                                                 // width_adapter_007:in_ready -> id_router_009:src_ready
	wire         width_adapter_007_src_endofpacket;                                                       // width_adapter_007:out_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         width_adapter_007_src_valid;                                                             // width_adapter_007:out_valid -> rsp_xbar_demux_009:sink_valid
	wire         width_adapter_007_src_startofpacket;                                                     // width_adapter_007:out_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [92:0] width_adapter_007_src_data;                                                              // width_adapter_007:out_data -> rsp_xbar_demux_009:sink_data
	wire         width_adapter_007_src_ready;                                                             // rsp_xbar_demux_009:sink_ready -> width_adapter_007:out_ready
	wire  [57:0] width_adapter_007_src_channel;                                                           // width_adapter_007:out_channel -> rsp_xbar_demux_009:sink_channel
	wire         cmd_xbar_demux_src10_ready;                                                              // width_adapter_008:in_ready -> cmd_xbar_demux:src10_ready
	wire         width_adapter_008_src_endofpacket;                                                       // width_adapter_008:out_endofpacket -> burst_adapter_011:sink0_endofpacket
	wire         width_adapter_008_src_valid;                                                             // width_adapter_008:out_valid -> burst_adapter_011:sink0_valid
	wire         width_adapter_008_src_startofpacket;                                                     // width_adapter_008:out_startofpacket -> burst_adapter_011:sink0_startofpacket
	wire  [65:0] width_adapter_008_src_data;                                                              // width_adapter_008:out_data -> burst_adapter_011:sink0_data
	wire         width_adapter_008_src_ready;                                                             // burst_adapter_011:sink0_ready -> width_adapter_008:out_ready
	wire  [57:0] width_adapter_008_src_channel;                                                           // width_adapter_008:out_channel -> burst_adapter_011:sink0_channel
	wire         id_router_010_src_endofpacket;                                                           // id_router_010:src_endofpacket -> width_adapter_009:in_endofpacket
	wire         id_router_010_src_valid;                                                                 // id_router_010:src_valid -> width_adapter_009:in_valid
	wire         id_router_010_src_startofpacket;                                                         // id_router_010:src_startofpacket -> width_adapter_009:in_startofpacket
	wire  [65:0] id_router_010_src_data;                                                                  // id_router_010:src_data -> width_adapter_009:in_data
	wire  [57:0] id_router_010_src_channel;                                                               // id_router_010:src_channel -> width_adapter_009:in_channel
	wire         id_router_010_src_ready;                                                                 // width_adapter_009:in_ready -> id_router_010:src_ready
	wire         width_adapter_009_src_endofpacket;                                                       // width_adapter_009:out_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         width_adapter_009_src_valid;                                                             // width_adapter_009:out_valid -> rsp_xbar_demux_010:sink_valid
	wire         width_adapter_009_src_startofpacket;                                                     // width_adapter_009:out_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [92:0] width_adapter_009_src_data;                                                              // width_adapter_009:out_data -> rsp_xbar_demux_010:sink_data
	wire         width_adapter_009_src_ready;                                                             // rsp_xbar_demux_010:sink_ready -> width_adapter_009:out_ready
	wire  [57:0] width_adapter_009_src_channel;                                                           // width_adapter_009:out_channel -> rsp_xbar_demux_010:sink_channel
	wire         cmd_xbar_demux_src11_ready;                                                              // width_adapter_010:in_ready -> cmd_xbar_demux:src11_ready
	wire         width_adapter_010_src_endofpacket;                                                       // width_adapter_010:out_endofpacket -> burst_adapter_049:sink0_endofpacket
	wire         width_adapter_010_src_valid;                                                             // width_adapter_010:out_valid -> burst_adapter_049:sink0_valid
	wire         width_adapter_010_src_startofpacket;                                                     // width_adapter_010:out_startofpacket -> burst_adapter_049:sink0_startofpacket
	wire  [65:0] width_adapter_010_src_data;                                                              // width_adapter_010:out_data -> burst_adapter_049:sink0_data
	wire         width_adapter_010_src_ready;                                                             // burst_adapter_049:sink0_ready -> width_adapter_010:out_ready
	wire  [57:0] width_adapter_010_src_channel;                                                           // width_adapter_010:out_channel -> burst_adapter_049:sink0_channel
	wire         id_router_011_src_endofpacket;                                                           // id_router_011:src_endofpacket -> width_adapter_011:in_endofpacket
	wire         id_router_011_src_valid;                                                                 // id_router_011:src_valid -> width_adapter_011:in_valid
	wire         id_router_011_src_startofpacket;                                                         // id_router_011:src_startofpacket -> width_adapter_011:in_startofpacket
	wire  [65:0] id_router_011_src_data;                                                                  // id_router_011:src_data -> width_adapter_011:in_data
	wire  [57:0] id_router_011_src_channel;                                                               // id_router_011:src_channel -> width_adapter_011:in_channel
	wire         id_router_011_src_ready;                                                                 // width_adapter_011:in_ready -> id_router_011:src_ready
	wire         width_adapter_011_src_endofpacket;                                                       // width_adapter_011:out_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         width_adapter_011_src_valid;                                                             // width_adapter_011:out_valid -> rsp_xbar_demux_011:sink_valid
	wire         width_adapter_011_src_startofpacket;                                                     // width_adapter_011:out_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [92:0] width_adapter_011_src_data;                                                              // width_adapter_011:out_data -> rsp_xbar_demux_011:sink_data
	wire         width_adapter_011_src_ready;                                                             // rsp_xbar_demux_011:sink_ready -> width_adapter_011:out_ready
	wire  [57:0] width_adapter_011_src_channel;                                                           // width_adapter_011:out_channel -> rsp_xbar_demux_011:sink_channel
	wire         cmd_xbar_demux_src12_ready;                                                              // width_adapter_012:in_ready -> cmd_xbar_demux:src12_ready
	wire         width_adapter_012_src_endofpacket;                                                       // width_adapter_012:out_endofpacket -> burst_adapter_010:sink0_endofpacket
	wire         width_adapter_012_src_valid;                                                             // width_adapter_012:out_valid -> burst_adapter_010:sink0_valid
	wire         width_adapter_012_src_startofpacket;                                                     // width_adapter_012:out_startofpacket -> burst_adapter_010:sink0_startofpacket
	wire  [65:0] width_adapter_012_src_data;                                                              // width_adapter_012:out_data -> burst_adapter_010:sink0_data
	wire         width_adapter_012_src_ready;                                                             // burst_adapter_010:sink0_ready -> width_adapter_012:out_ready
	wire  [57:0] width_adapter_012_src_channel;                                                           // width_adapter_012:out_channel -> burst_adapter_010:sink0_channel
	wire         id_router_012_src_endofpacket;                                                           // id_router_012:src_endofpacket -> width_adapter_013:in_endofpacket
	wire         id_router_012_src_valid;                                                                 // id_router_012:src_valid -> width_adapter_013:in_valid
	wire         id_router_012_src_startofpacket;                                                         // id_router_012:src_startofpacket -> width_adapter_013:in_startofpacket
	wire  [65:0] id_router_012_src_data;                                                                  // id_router_012:src_data -> width_adapter_013:in_data
	wire  [57:0] id_router_012_src_channel;                                                               // id_router_012:src_channel -> width_adapter_013:in_channel
	wire         id_router_012_src_ready;                                                                 // width_adapter_013:in_ready -> id_router_012:src_ready
	wire         width_adapter_013_src_endofpacket;                                                       // width_adapter_013:out_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         width_adapter_013_src_valid;                                                             // width_adapter_013:out_valid -> rsp_xbar_demux_012:sink_valid
	wire         width_adapter_013_src_startofpacket;                                                     // width_adapter_013:out_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [92:0] width_adapter_013_src_data;                                                              // width_adapter_013:out_data -> rsp_xbar_demux_012:sink_data
	wire         width_adapter_013_src_ready;                                                             // rsp_xbar_demux_012:sink_ready -> width_adapter_013:out_ready
	wire  [57:0] width_adapter_013_src_channel;                                                           // width_adapter_013:out_channel -> rsp_xbar_demux_012:sink_channel
	wire         cmd_xbar_demux_src13_ready;                                                              // width_adapter_014:in_ready -> cmd_xbar_demux:src13_ready
	wire         width_adapter_014_src_endofpacket;                                                       // width_adapter_014:out_endofpacket -> burst_adapter_023:sink0_endofpacket
	wire         width_adapter_014_src_valid;                                                             // width_adapter_014:out_valid -> burst_adapter_023:sink0_valid
	wire         width_adapter_014_src_startofpacket;                                                     // width_adapter_014:out_startofpacket -> burst_adapter_023:sink0_startofpacket
	wire  [65:0] width_adapter_014_src_data;                                                              // width_adapter_014:out_data -> burst_adapter_023:sink0_data
	wire         width_adapter_014_src_ready;                                                             // burst_adapter_023:sink0_ready -> width_adapter_014:out_ready
	wire  [57:0] width_adapter_014_src_channel;                                                           // width_adapter_014:out_channel -> burst_adapter_023:sink0_channel
	wire         id_router_013_src_endofpacket;                                                           // id_router_013:src_endofpacket -> width_adapter_015:in_endofpacket
	wire         id_router_013_src_valid;                                                                 // id_router_013:src_valid -> width_adapter_015:in_valid
	wire         id_router_013_src_startofpacket;                                                         // id_router_013:src_startofpacket -> width_adapter_015:in_startofpacket
	wire  [65:0] id_router_013_src_data;                                                                  // id_router_013:src_data -> width_adapter_015:in_data
	wire  [57:0] id_router_013_src_channel;                                                               // id_router_013:src_channel -> width_adapter_015:in_channel
	wire         id_router_013_src_ready;                                                                 // width_adapter_015:in_ready -> id_router_013:src_ready
	wire         width_adapter_015_src_endofpacket;                                                       // width_adapter_015:out_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         width_adapter_015_src_valid;                                                             // width_adapter_015:out_valid -> rsp_xbar_demux_013:sink_valid
	wire         width_adapter_015_src_startofpacket;                                                     // width_adapter_015:out_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [92:0] width_adapter_015_src_data;                                                              // width_adapter_015:out_data -> rsp_xbar_demux_013:sink_data
	wire         width_adapter_015_src_ready;                                                             // rsp_xbar_demux_013:sink_ready -> width_adapter_015:out_ready
	wire  [57:0] width_adapter_015_src_channel;                                                           // width_adapter_015:out_channel -> rsp_xbar_demux_013:sink_channel
	wire         cmd_xbar_demux_src14_ready;                                                              // width_adapter_016:in_ready -> cmd_xbar_demux:src14_ready
	wire         width_adapter_016_src_endofpacket;                                                       // width_adapter_016:out_endofpacket -> burst_adapter_043:sink0_endofpacket
	wire         width_adapter_016_src_valid;                                                             // width_adapter_016:out_valid -> burst_adapter_043:sink0_valid
	wire         width_adapter_016_src_startofpacket;                                                     // width_adapter_016:out_startofpacket -> burst_adapter_043:sink0_startofpacket
	wire  [65:0] width_adapter_016_src_data;                                                              // width_adapter_016:out_data -> burst_adapter_043:sink0_data
	wire         width_adapter_016_src_ready;                                                             // burst_adapter_043:sink0_ready -> width_adapter_016:out_ready
	wire  [57:0] width_adapter_016_src_channel;                                                           // width_adapter_016:out_channel -> burst_adapter_043:sink0_channel
	wire         id_router_014_src_endofpacket;                                                           // id_router_014:src_endofpacket -> width_adapter_017:in_endofpacket
	wire         id_router_014_src_valid;                                                                 // id_router_014:src_valid -> width_adapter_017:in_valid
	wire         id_router_014_src_startofpacket;                                                         // id_router_014:src_startofpacket -> width_adapter_017:in_startofpacket
	wire  [65:0] id_router_014_src_data;                                                                  // id_router_014:src_data -> width_adapter_017:in_data
	wire  [57:0] id_router_014_src_channel;                                                               // id_router_014:src_channel -> width_adapter_017:in_channel
	wire         id_router_014_src_ready;                                                                 // width_adapter_017:in_ready -> id_router_014:src_ready
	wire         width_adapter_017_src_endofpacket;                                                       // width_adapter_017:out_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire         width_adapter_017_src_valid;                                                             // width_adapter_017:out_valid -> rsp_xbar_demux_014:sink_valid
	wire         width_adapter_017_src_startofpacket;                                                     // width_adapter_017:out_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [92:0] width_adapter_017_src_data;                                                              // width_adapter_017:out_data -> rsp_xbar_demux_014:sink_data
	wire         width_adapter_017_src_ready;                                                             // rsp_xbar_demux_014:sink_ready -> width_adapter_017:out_ready
	wire  [57:0] width_adapter_017_src_channel;                                                           // width_adapter_017:out_channel -> rsp_xbar_demux_014:sink_channel
	wire         cmd_xbar_demux_src15_ready;                                                              // width_adapter_018:in_ready -> cmd_xbar_demux:src15_ready
	wire         width_adapter_018_src_endofpacket;                                                       // width_adapter_018:out_endofpacket -> burst_adapter_042:sink0_endofpacket
	wire         width_adapter_018_src_valid;                                                             // width_adapter_018:out_valid -> burst_adapter_042:sink0_valid
	wire         width_adapter_018_src_startofpacket;                                                     // width_adapter_018:out_startofpacket -> burst_adapter_042:sink0_startofpacket
	wire  [65:0] width_adapter_018_src_data;                                                              // width_adapter_018:out_data -> burst_adapter_042:sink0_data
	wire         width_adapter_018_src_ready;                                                             // burst_adapter_042:sink0_ready -> width_adapter_018:out_ready
	wire  [57:0] width_adapter_018_src_channel;                                                           // width_adapter_018:out_channel -> burst_adapter_042:sink0_channel
	wire         id_router_015_src_endofpacket;                                                           // id_router_015:src_endofpacket -> width_adapter_019:in_endofpacket
	wire         id_router_015_src_valid;                                                                 // id_router_015:src_valid -> width_adapter_019:in_valid
	wire         id_router_015_src_startofpacket;                                                         // id_router_015:src_startofpacket -> width_adapter_019:in_startofpacket
	wire  [65:0] id_router_015_src_data;                                                                  // id_router_015:src_data -> width_adapter_019:in_data
	wire  [57:0] id_router_015_src_channel;                                                               // id_router_015:src_channel -> width_adapter_019:in_channel
	wire         id_router_015_src_ready;                                                                 // width_adapter_019:in_ready -> id_router_015:src_ready
	wire         width_adapter_019_src_endofpacket;                                                       // width_adapter_019:out_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire         width_adapter_019_src_valid;                                                             // width_adapter_019:out_valid -> rsp_xbar_demux_015:sink_valid
	wire         width_adapter_019_src_startofpacket;                                                     // width_adapter_019:out_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [92:0] width_adapter_019_src_data;                                                              // width_adapter_019:out_data -> rsp_xbar_demux_015:sink_data
	wire         width_adapter_019_src_ready;                                                             // rsp_xbar_demux_015:sink_ready -> width_adapter_019:out_ready
	wire  [57:0] width_adapter_019_src_channel;                                                           // width_adapter_019:out_channel -> rsp_xbar_demux_015:sink_channel
	wire         cmd_xbar_demux_src16_ready;                                                              // width_adapter_020:in_ready -> cmd_xbar_demux:src16_ready
	wire         width_adapter_020_src_endofpacket;                                                       // width_adapter_020:out_endofpacket -> burst_adapter_007:sink0_endofpacket
	wire         width_adapter_020_src_valid;                                                             // width_adapter_020:out_valid -> burst_adapter_007:sink0_valid
	wire         width_adapter_020_src_startofpacket;                                                     // width_adapter_020:out_startofpacket -> burst_adapter_007:sink0_startofpacket
	wire  [65:0] width_adapter_020_src_data;                                                              // width_adapter_020:out_data -> burst_adapter_007:sink0_data
	wire         width_adapter_020_src_ready;                                                             // burst_adapter_007:sink0_ready -> width_adapter_020:out_ready
	wire  [57:0] width_adapter_020_src_channel;                                                           // width_adapter_020:out_channel -> burst_adapter_007:sink0_channel
	wire         id_router_016_src_endofpacket;                                                           // id_router_016:src_endofpacket -> width_adapter_021:in_endofpacket
	wire         id_router_016_src_valid;                                                                 // id_router_016:src_valid -> width_adapter_021:in_valid
	wire         id_router_016_src_startofpacket;                                                         // id_router_016:src_startofpacket -> width_adapter_021:in_startofpacket
	wire  [65:0] id_router_016_src_data;                                                                  // id_router_016:src_data -> width_adapter_021:in_data
	wire  [57:0] id_router_016_src_channel;                                                               // id_router_016:src_channel -> width_adapter_021:in_channel
	wire         id_router_016_src_ready;                                                                 // width_adapter_021:in_ready -> id_router_016:src_ready
	wire         width_adapter_021_src_endofpacket;                                                       // width_adapter_021:out_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire         width_adapter_021_src_valid;                                                             // width_adapter_021:out_valid -> rsp_xbar_demux_016:sink_valid
	wire         width_adapter_021_src_startofpacket;                                                     // width_adapter_021:out_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [92:0] width_adapter_021_src_data;                                                              // width_adapter_021:out_data -> rsp_xbar_demux_016:sink_data
	wire         width_adapter_021_src_ready;                                                             // rsp_xbar_demux_016:sink_ready -> width_adapter_021:out_ready
	wire  [57:0] width_adapter_021_src_channel;                                                           // width_adapter_021:out_channel -> rsp_xbar_demux_016:sink_channel
	wire         cmd_xbar_demux_src17_ready;                                                              // width_adapter_022:in_ready -> cmd_xbar_demux:src17_ready
	wire         width_adapter_022_src_endofpacket;                                                       // width_adapter_022:out_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire         width_adapter_022_src_valid;                                                             // width_adapter_022:out_valid -> burst_adapter_003:sink0_valid
	wire         width_adapter_022_src_startofpacket;                                                     // width_adapter_022:out_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire  [65:0] width_adapter_022_src_data;                                                              // width_adapter_022:out_data -> burst_adapter_003:sink0_data
	wire         width_adapter_022_src_ready;                                                             // burst_adapter_003:sink0_ready -> width_adapter_022:out_ready
	wire  [57:0] width_adapter_022_src_channel;                                                           // width_adapter_022:out_channel -> burst_adapter_003:sink0_channel
	wire         id_router_017_src_endofpacket;                                                           // id_router_017:src_endofpacket -> width_adapter_023:in_endofpacket
	wire         id_router_017_src_valid;                                                                 // id_router_017:src_valid -> width_adapter_023:in_valid
	wire         id_router_017_src_startofpacket;                                                         // id_router_017:src_startofpacket -> width_adapter_023:in_startofpacket
	wire  [65:0] id_router_017_src_data;                                                                  // id_router_017:src_data -> width_adapter_023:in_data
	wire  [57:0] id_router_017_src_channel;                                                               // id_router_017:src_channel -> width_adapter_023:in_channel
	wire         id_router_017_src_ready;                                                                 // width_adapter_023:in_ready -> id_router_017:src_ready
	wire         width_adapter_023_src_endofpacket;                                                       // width_adapter_023:out_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire         width_adapter_023_src_valid;                                                             // width_adapter_023:out_valid -> rsp_xbar_demux_017:sink_valid
	wire         width_adapter_023_src_startofpacket;                                                     // width_adapter_023:out_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [92:0] width_adapter_023_src_data;                                                              // width_adapter_023:out_data -> rsp_xbar_demux_017:sink_data
	wire         width_adapter_023_src_ready;                                                             // rsp_xbar_demux_017:sink_ready -> width_adapter_023:out_ready
	wire  [57:0] width_adapter_023_src_channel;                                                           // width_adapter_023:out_channel -> rsp_xbar_demux_017:sink_channel
	wire         cmd_xbar_demux_src18_ready;                                                              // width_adapter_024:in_ready -> cmd_xbar_demux:src18_ready
	wire         width_adapter_024_src_endofpacket;                                                       // width_adapter_024:out_endofpacket -> burst_adapter_046:sink0_endofpacket
	wire         width_adapter_024_src_valid;                                                             // width_adapter_024:out_valid -> burst_adapter_046:sink0_valid
	wire         width_adapter_024_src_startofpacket;                                                     // width_adapter_024:out_startofpacket -> burst_adapter_046:sink0_startofpacket
	wire  [65:0] width_adapter_024_src_data;                                                              // width_adapter_024:out_data -> burst_adapter_046:sink0_data
	wire         width_adapter_024_src_ready;                                                             // burst_adapter_046:sink0_ready -> width_adapter_024:out_ready
	wire  [57:0] width_adapter_024_src_channel;                                                           // width_adapter_024:out_channel -> burst_adapter_046:sink0_channel
	wire         id_router_018_src_endofpacket;                                                           // id_router_018:src_endofpacket -> width_adapter_025:in_endofpacket
	wire         id_router_018_src_valid;                                                                 // id_router_018:src_valid -> width_adapter_025:in_valid
	wire         id_router_018_src_startofpacket;                                                         // id_router_018:src_startofpacket -> width_adapter_025:in_startofpacket
	wire  [65:0] id_router_018_src_data;                                                                  // id_router_018:src_data -> width_adapter_025:in_data
	wire  [57:0] id_router_018_src_channel;                                                               // id_router_018:src_channel -> width_adapter_025:in_channel
	wire         id_router_018_src_ready;                                                                 // width_adapter_025:in_ready -> id_router_018:src_ready
	wire         width_adapter_025_src_endofpacket;                                                       // width_adapter_025:out_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire         width_adapter_025_src_valid;                                                             // width_adapter_025:out_valid -> rsp_xbar_demux_018:sink_valid
	wire         width_adapter_025_src_startofpacket;                                                     // width_adapter_025:out_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [92:0] width_adapter_025_src_data;                                                              // width_adapter_025:out_data -> rsp_xbar_demux_018:sink_data
	wire         width_adapter_025_src_ready;                                                             // rsp_xbar_demux_018:sink_ready -> width_adapter_025:out_ready
	wire  [57:0] width_adapter_025_src_channel;                                                           // width_adapter_025:out_channel -> rsp_xbar_demux_018:sink_channel
	wire         cmd_xbar_demux_src19_ready;                                                              // width_adapter_026:in_ready -> cmd_xbar_demux:src19_ready
	wire         width_adapter_026_src_endofpacket;                                                       // width_adapter_026:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire         width_adapter_026_src_valid;                                                             // width_adapter_026:out_valid -> burst_adapter_002:sink0_valid
	wire         width_adapter_026_src_startofpacket;                                                     // width_adapter_026:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire  [65:0] width_adapter_026_src_data;                                                              // width_adapter_026:out_data -> burst_adapter_002:sink0_data
	wire         width_adapter_026_src_ready;                                                             // burst_adapter_002:sink0_ready -> width_adapter_026:out_ready
	wire  [57:0] width_adapter_026_src_channel;                                                           // width_adapter_026:out_channel -> burst_adapter_002:sink0_channel
	wire         id_router_019_src_endofpacket;                                                           // id_router_019:src_endofpacket -> width_adapter_027:in_endofpacket
	wire         id_router_019_src_valid;                                                                 // id_router_019:src_valid -> width_adapter_027:in_valid
	wire         id_router_019_src_startofpacket;                                                         // id_router_019:src_startofpacket -> width_adapter_027:in_startofpacket
	wire  [65:0] id_router_019_src_data;                                                                  // id_router_019:src_data -> width_adapter_027:in_data
	wire  [57:0] id_router_019_src_channel;                                                               // id_router_019:src_channel -> width_adapter_027:in_channel
	wire         id_router_019_src_ready;                                                                 // width_adapter_027:in_ready -> id_router_019:src_ready
	wire         width_adapter_027_src_endofpacket;                                                       // width_adapter_027:out_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire         width_adapter_027_src_valid;                                                             // width_adapter_027:out_valid -> rsp_xbar_demux_019:sink_valid
	wire         width_adapter_027_src_startofpacket;                                                     // width_adapter_027:out_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [92:0] width_adapter_027_src_data;                                                              // width_adapter_027:out_data -> rsp_xbar_demux_019:sink_data
	wire         width_adapter_027_src_ready;                                                             // rsp_xbar_demux_019:sink_ready -> width_adapter_027:out_ready
	wire  [57:0] width_adapter_027_src_channel;                                                           // width_adapter_027:out_channel -> rsp_xbar_demux_019:sink_channel
	wire         cmd_xbar_demux_src20_ready;                                                              // width_adapter_028:in_ready -> cmd_xbar_demux:src20_ready
	wire         width_adapter_028_src_endofpacket;                                                       // width_adapter_028:out_endofpacket -> burst_adapter_027:sink0_endofpacket
	wire         width_adapter_028_src_valid;                                                             // width_adapter_028:out_valid -> burst_adapter_027:sink0_valid
	wire         width_adapter_028_src_startofpacket;                                                     // width_adapter_028:out_startofpacket -> burst_adapter_027:sink0_startofpacket
	wire  [65:0] width_adapter_028_src_data;                                                              // width_adapter_028:out_data -> burst_adapter_027:sink0_data
	wire         width_adapter_028_src_ready;                                                             // burst_adapter_027:sink0_ready -> width_adapter_028:out_ready
	wire  [57:0] width_adapter_028_src_channel;                                                           // width_adapter_028:out_channel -> burst_adapter_027:sink0_channel
	wire         id_router_020_src_endofpacket;                                                           // id_router_020:src_endofpacket -> width_adapter_029:in_endofpacket
	wire         id_router_020_src_valid;                                                                 // id_router_020:src_valid -> width_adapter_029:in_valid
	wire         id_router_020_src_startofpacket;                                                         // id_router_020:src_startofpacket -> width_adapter_029:in_startofpacket
	wire  [65:0] id_router_020_src_data;                                                                  // id_router_020:src_data -> width_adapter_029:in_data
	wire  [57:0] id_router_020_src_channel;                                                               // id_router_020:src_channel -> width_adapter_029:in_channel
	wire         id_router_020_src_ready;                                                                 // width_adapter_029:in_ready -> id_router_020:src_ready
	wire         width_adapter_029_src_endofpacket;                                                       // width_adapter_029:out_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire         width_adapter_029_src_valid;                                                             // width_adapter_029:out_valid -> rsp_xbar_demux_020:sink_valid
	wire         width_adapter_029_src_startofpacket;                                                     // width_adapter_029:out_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [92:0] width_adapter_029_src_data;                                                              // width_adapter_029:out_data -> rsp_xbar_demux_020:sink_data
	wire         width_adapter_029_src_ready;                                                             // rsp_xbar_demux_020:sink_ready -> width_adapter_029:out_ready
	wire  [57:0] width_adapter_029_src_channel;                                                           // width_adapter_029:out_channel -> rsp_xbar_demux_020:sink_channel
	wire         cmd_xbar_demux_src21_ready;                                                              // width_adapter_030:in_ready -> cmd_xbar_demux:src21_ready
	wire         width_adapter_030_src_endofpacket;                                                       // width_adapter_030:out_endofpacket -> burst_adapter_040:sink0_endofpacket
	wire         width_adapter_030_src_valid;                                                             // width_adapter_030:out_valid -> burst_adapter_040:sink0_valid
	wire         width_adapter_030_src_startofpacket;                                                     // width_adapter_030:out_startofpacket -> burst_adapter_040:sink0_startofpacket
	wire  [65:0] width_adapter_030_src_data;                                                              // width_adapter_030:out_data -> burst_adapter_040:sink0_data
	wire         width_adapter_030_src_ready;                                                             // burst_adapter_040:sink0_ready -> width_adapter_030:out_ready
	wire  [57:0] width_adapter_030_src_channel;                                                           // width_adapter_030:out_channel -> burst_adapter_040:sink0_channel
	wire         id_router_021_src_endofpacket;                                                           // id_router_021:src_endofpacket -> width_adapter_031:in_endofpacket
	wire         id_router_021_src_valid;                                                                 // id_router_021:src_valid -> width_adapter_031:in_valid
	wire         id_router_021_src_startofpacket;                                                         // id_router_021:src_startofpacket -> width_adapter_031:in_startofpacket
	wire  [65:0] id_router_021_src_data;                                                                  // id_router_021:src_data -> width_adapter_031:in_data
	wire  [57:0] id_router_021_src_channel;                                                               // id_router_021:src_channel -> width_adapter_031:in_channel
	wire         id_router_021_src_ready;                                                                 // width_adapter_031:in_ready -> id_router_021:src_ready
	wire         width_adapter_031_src_endofpacket;                                                       // width_adapter_031:out_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire         width_adapter_031_src_valid;                                                             // width_adapter_031:out_valid -> rsp_xbar_demux_021:sink_valid
	wire         width_adapter_031_src_startofpacket;                                                     // width_adapter_031:out_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [92:0] width_adapter_031_src_data;                                                              // width_adapter_031:out_data -> rsp_xbar_demux_021:sink_data
	wire         width_adapter_031_src_ready;                                                             // rsp_xbar_demux_021:sink_ready -> width_adapter_031:out_ready
	wire  [57:0] width_adapter_031_src_channel;                                                           // width_adapter_031:out_channel -> rsp_xbar_demux_021:sink_channel
	wire         cmd_xbar_demux_src22_ready;                                                              // width_adapter_032:in_ready -> cmd_xbar_demux:src22_ready
	wire         width_adapter_032_src_endofpacket;                                                       // width_adapter_032:out_endofpacket -> burst_adapter_014:sink0_endofpacket
	wire         width_adapter_032_src_valid;                                                             // width_adapter_032:out_valid -> burst_adapter_014:sink0_valid
	wire         width_adapter_032_src_startofpacket;                                                     // width_adapter_032:out_startofpacket -> burst_adapter_014:sink0_startofpacket
	wire  [65:0] width_adapter_032_src_data;                                                              // width_adapter_032:out_data -> burst_adapter_014:sink0_data
	wire         width_adapter_032_src_ready;                                                             // burst_adapter_014:sink0_ready -> width_adapter_032:out_ready
	wire  [57:0] width_adapter_032_src_channel;                                                           // width_adapter_032:out_channel -> burst_adapter_014:sink0_channel
	wire         id_router_022_src_endofpacket;                                                           // id_router_022:src_endofpacket -> width_adapter_033:in_endofpacket
	wire         id_router_022_src_valid;                                                                 // id_router_022:src_valid -> width_adapter_033:in_valid
	wire         id_router_022_src_startofpacket;                                                         // id_router_022:src_startofpacket -> width_adapter_033:in_startofpacket
	wire  [65:0] id_router_022_src_data;                                                                  // id_router_022:src_data -> width_adapter_033:in_data
	wire  [57:0] id_router_022_src_channel;                                                               // id_router_022:src_channel -> width_adapter_033:in_channel
	wire         id_router_022_src_ready;                                                                 // width_adapter_033:in_ready -> id_router_022:src_ready
	wire         width_adapter_033_src_endofpacket;                                                       // width_adapter_033:out_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire         width_adapter_033_src_valid;                                                             // width_adapter_033:out_valid -> rsp_xbar_demux_022:sink_valid
	wire         width_adapter_033_src_startofpacket;                                                     // width_adapter_033:out_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [92:0] width_adapter_033_src_data;                                                              // width_adapter_033:out_data -> rsp_xbar_demux_022:sink_data
	wire         width_adapter_033_src_ready;                                                             // rsp_xbar_demux_022:sink_ready -> width_adapter_033:out_ready
	wire  [57:0] width_adapter_033_src_channel;                                                           // width_adapter_033:out_channel -> rsp_xbar_demux_022:sink_channel
	wire         cmd_xbar_demux_src23_ready;                                                              // width_adapter_034:in_ready -> cmd_xbar_demux:src23_ready
	wire         width_adapter_034_src_endofpacket;                                                       // width_adapter_034:out_endofpacket -> burst_adapter_047:sink0_endofpacket
	wire         width_adapter_034_src_valid;                                                             // width_adapter_034:out_valid -> burst_adapter_047:sink0_valid
	wire         width_adapter_034_src_startofpacket;                                                     // width_adapter_034:out_startofpacket -> burst_adapter_047:sink0_startofpacket
	wire  [65:0] width_adapter_034_src_data;                                                              // width_adapter_034:out_data -> burst_adapter_047:sink0_data
	wire         width_adapter_034_src_ready;                                                             // burst_adapter_047:sink0_ready -> width_adapter_034:out_ready
	wire  [57:0] width_adapter_034_src_channel;                                                           // width_adapter_034:out_channel -> burst_adapter_047:sink0_channel
	wire         id_router_023_src_endofpacket;                                                           // id_router_023:src_endofpacket -> width_adapter_035:in_endofpacket
	wire         id_router_023_src_valid;                                                                 // id_router_023:src_valid -> width_adapter_035:in_valid
	wire         id_router_023_src_startofpacket;                                                         // id_router_023:src_startofpacket -> width_adapter_035:in_startofpacket
	wire  [65:0] id_router_023_src_data;                                                                  // id_router_023:src_data -> width_adapter_035:in_data
	wire  [57:0] id_router_023_src_channel;                                                               // id_router_023:src_channel -> width_adapter_035:in_channel
	wire         id_router_023_src_ready;                                                                 // width_adapter_035:in_ready -> id_router_023:src_ready
	wire         width_adapter_035_src_endofpacket;                                                       // width_adapter_035:out_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire         width_adapter_035_src_valid;                                                             // width_adapter_035:out_valid -> rsp_xbar_demux_023:sink_valid
	wire         width_adapter_035_src_startofpacket;                                                     // width_adapter_035:out_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire  [92:0] width_adapter_035_src_data;                                                              // width_adapter_035:out_data -> rsp_xbar_demux_023:sink_data
	wire         width_adapter_035_src_ready;                                                             // rsp_xbar_demux_023:sink_ready -> width_adapter_035:out_ready
	wire  [57:0] width_adapter_035_src_channel;                                                           // width_adapter_035:out_channel -> rsp_xbar_demux_023:sink_channel
	wire         cmd_xbar_demux_src24_ready;                                                              // width_adapter_036:in_ready -> cmd_xbar_demux:src24_ready
	wire         width_adapter_036_src_endofpacket;                                                       // width_adapter_036:out_endofpacket -> burst_adapter_051:sink0_endofpacket
	wire         width_adapter_036_src_valid;                                                             // width_adapter_036:out_valid -> burst_adapter_051:sink0_valid
	wire         width_adapter_036_src_startofpacket;                                                     // width_adapter_036:out_startofpacket -> burst_adapter_051:sink0_startofpacket
	wire  [65:0] width_adapter_036_src_data;                                                              // width_adapter_036:out_data -> burst_adapter_051:sink0_data
	wire         width_adapter_036_src_ready;                                                             // burst_adapter_051:sink0_ready -> width_adapter_036:out_ready
	wire  [57:0] width_adapter_036_src_channel;                                                           // width_adapter_036:out_channel -> burst_adapter_051:sink0_channel
	wire         id_router_024_src_endofpacket;                                                           // id_router_024:src_endofpacket -> width_adapter_037:in_endofpacket
	wire         id_router_024_src_valid;                                                                 // id_router_024:src_valid -> width_adapter_037:in_valid
	wire         id_router_024_src_startofpacket;                                                         // id_router_024:src_startofpacket -> width_adapter_037:in_startofpacket
	wire  [65:0] id_router_024_src_data;                                                                  // id_router_024:src_data -> width_adapter_037:in_data
	wire  [57:0] id_router_024_src_channel;                                                               // id_router_024:src_channel -> width_adapter_037:in_channel
	wire         id_router_024_src_ready;                                                                 // width_adapter_037:in_ready -> id_router_024:src_ready
	wire         width_adapter_037_src_endofpacket;                                                       // width_adapter_037:out_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire         width_adapter_037_src_valid;                                                             // width_adapter_037:out_valid -> rsp_xbar_demux_024:sink_valid
	wire         width_adapter_037_src_startofpacket;                                                     // width_adapter_037:out_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire  [92:0] width_adapter_037_src_data;                                                              // width_adapter_037:out_data -> rsp_xbar_demux_024:sink_data
	wire         width_adapter_037_src_ready;                                                             // rsp_xbar_demux_024:sink_ready -> width_adapter_037:out_ready
	wire  [57:0] width_adapter_037_src_channel;                                                           // width_adapter_037:out_channel -> rsp_xbar_demux_024:sink_channel
	wire         cmd_xbar_demux_src25_ready;                                                              // width_adapter_038:in_ready -> cmd_xbar_demux:src25_ready
	wire         width_adapter_038_src_endofpacket;                                                       // width_adapter_038:out_endofpacket -> burst_adapter_008:sink0_endofpacket
	wire         width_adapter_038_src_valid;                                                             // width_adapter_038:out_valid -> burst_adapter_008:sink0_valid
	wire         width_adapter_038_src_startofpacket;                                                     // width_adapter_038:out_startofpacket -> burst_adapter_008:sink0_startofpacket
	wire  [65:0] width_adapter_038_src_data;                                                              // width_adapter_038:out_data -> burst_adapter_008:sink0_data
	wire         width_adapter_038_src_ready;                                                             // burst_adapter_008:sink0_ready -> width_adapter_038:out_ready
	wire  [57:0] width_adapter_038_src_channel;                                                           // width_adapter_038:out_channel -> burst_adapter_008:sink0_channel
	wire         id_router_025_src_endofpacket;                                                           // id_router_025:src_endofpacket -> width_adapter_039:in_endofpacket
	wire         id_router_025_src_valid;                                                                 // id_router_025:src_valid -> width_adapter_039:in_valid
	wire         id_router_025_src_startofpacket;                                                         // id_router_025:src_startofpacket -> width_adapter_039:in_startofpacket
	wire  [65:0] id_router_025_src_data;                                                                  // id_router_025:src_data -> width_adapter_039:in_data
	wire  [57:0] id_router_025_src_channel;                                                               // id_router_025:src_channel -> width_adapter_039:in_channel
	wire         id_router_025_src_ready;                                                                 // width_adapter_039:in_ready -> id_router_025:src_ready
	wire         width_adapter_039_src_endofpacket;                                                       // width_adapter_039:out_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire         width_adapter_039_src_valid;                                                             // width_adapter_039:out_valid -> rsp_xbar_demux_025:sink_valid
	wire         width_adapter_039_src_startofpacket;                                                     // width_adapter_039:out_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire  [92:0] width_adapter_039_src_data;                                                              // width_adapter_039:out_data -> rsp_xbar_demux_025:sink_data
	wire         width_adapter_039_src_ready;                                                             // rsp_xbar_demux_025:sink_ready -> width_adapter_039:out_ready
	wire  [57:0] width_adapter_039_src_channel;                                                           // width_adapter_039:out_channel -> rsp_xbar_demux_025:sink_channel
	wire         cmd_xbar_demux_src26_ready;                                                              // width_adapter_040:in_ready -> cmd_xbar_demux:src26_ready
	wire         width_adapter_040_src_endofpacket;                                                       // width_adapter_040:out_endofpacket -> burst_adapter_012:sink0_endofpacket
	wire         width_adapter_040_src_valid;                                                             // width_adapter_040:out_valid -> burst_adapter_012:sink0_valid
	wire         width_adapter_040_src_startofpacket;                                                     // width_adapter_040:out_startofpacket -> burst_adapter_012:sink0_startofpacket
	wire  [65:0] width_adapter_040_src_data;                                                              // width_adapter_040:out_data -> burst_adapter_012:sink0_data
	wire         width_adapter_040_src_ready;                                                             // burst_adapter_012:sink0_ready -> width_adapter_040:out_ready
	wire  [57:0] width_adapter_040_src_channel;                                                           // width_adapter_040:out_channel -> burst_adapter_012:sink0_channel
	wire         id_router_026_src_endofpacket;                                                           // id_router_026:src_endofpacket -> width_adapter_041:in_endofpacket
	wire         id_router_026_src_valid;                                                                 // id_router_026:src_valid -> width_adapter_041:in_valid
	wire         id_router_026_src_startofpacket;                                                         // id_router_026:src_startofpacket -> width_adapter_041:in_startofpacket
	wire  [65:0] id_router_026_src_data;                                                                  // id_router_026:src_data -> width_adapter_041:in_data
	wire  [57:0] id_router_026_src_channel;                                                               // id_router_026:src_channel -> width_adapter_041:in_channel
	wire         id_router_026_src_ready;                                                                 // width_adapter_041:in_ready -> id_router_026:src_ready
	wire         width_adapter_041_src_endofpacket;                                                       // width_adapter_041:out_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	wire         width_adapter_041_src_valid;                                                             // width_adapter_041:out_valid -> rsp_xbar_demux_026:sink_valid
	wire         width_adapter_041_src_startofpacket;                                                     // width_adapter_041:out_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	wire  [92:0] width_adapter_041_src_data;                                                              // width_adapter_041:out_data -> rsp_xbar_demux_026:sink_data
	wire         width_adapter_041_src_ready;                                                             // rsp_xbar_demux_026:sink_ready -> width_adapter_041:out_ready
	wire  [57:0] width_adapter_041_src_channel;                                                           // width_adapter_041:out_channel -> rsp_xbar_demux_026:sink_channel
	wire         cmd_xbar_demux_src27_ready;                                                              // width_adapter_042:in_ready -> cmd_xbar_demux:src27_ready
	wire         width_adapter_042_src_endofpacket;                                                       // width_adapter_042:out_endofpacket -> burst_adapter_037:sink0_endofpacket
	wire         width_adapter_042_src_valid;                                                             // width_adapter_042:out_valid -> burst_adapter_037:sink0_valid
	wire         width_adapter_042_src_startofpacket;                                                     // width_adapter_042:out_startofpacket -> burst_adapter_037:sink0_startofpacket
	wire  [65:0] width_adapter_042_src_data;                                                              // width_adapter_042:out_data -> burst_adapter_037:sink0_data
	wire         width_adapter_042_src_ready;                                                             // burst_adapter_037:sink0_ready -> width_adapter_042:out_ready
	wire  [57:0] width_adapter_042_src_channel;                                                           // width_adapter_042:out_channel -> burst_adapter_037:sink0_channel
	wire         id_router_027_src_endofpacket;                                                           // id_router_027:src_endofpacket -> width_adapter_043:in_endofpacket
	wire         id_router_027_src_valid;                                                                 // id_router_027:src_valid -> width_adapter_043:in_valid
	wire         id_router_027_src_startofpacket;                                                         // id_router_027:src_startofpacket -> width_adapter_043:in_startofpacket
	wire  [65:0] id_router_027_src_data;                                                                  // id_router_027:src_data -> width_adapter_043:in_data
	wire  [57:0] id_router_027_src_channel;                                                               // id_router_027:src_channel -> width_adapter_043:in_channel
	wire         id_router_027_src_ready;                                                                 // width_adapter_043:in_ready -> id_router_027:src_ready
	wire         width_adapter_043_src_endofpacket;                                                       // width_adapter_043:out_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	wire         width_adapter_043_src_valid;                                                             // width_adapter_043:out_valid -> rsp_xbar_demux_027:sink_valid
	wire         width_adapter_043_src_startofpacket;                                                     // width_adapter_043:out_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	wire  [92:0] width_adapter_043_src_data;                                                              // width_adapter_043:out_data -> rsp_xbar_demux_027:sink_data
	wire         width_adapter_043_src_ready;                                                             // rsp_xbar_demux_027:sink_ready -> width_adapter_043:out_ready
	wire  [57:0] width_adapter_043_src_channel;                                                           // width_adapter_043:out_channel -> rsp_xbar_demux_027:sink_channel
	wire         cmd_xbar_demux_src28_ready;                                                              // width_adapter_044:in_ready -> cmd_xbar_demux:src28_ready
	wire         width_adapter_044_src_endofpacket;                                                       // width_adapter_044:out_endofpacket -> burst_adapter_033:sink0_endofpacket
	wire         width_adapter_044_src_valid;                                                             // width_adapter_044:out_valid -> burst_adapter_033:sink0_valid
	wire         width_adapter_044_src_startofpacket;                                                     // width_adapter_044:out_startofpacket -> burst_adapter_033:sink0_startofpacket
	wire  [65:0] width_adapter_044_src_data;                                                              // width_adapter_044:out_data -> burst_adapter_033:sink0_data
	wire         width_adapter_044_src_ready;                                                             // burst_adapter_033:sink0_ready -> width_adapter_044:out_ready
	wire  [57:0] width_adapter_044_src_channel;                                                           // width_adapter_044:out_channel -> burst_adapter_033:sink0_channel
	wire         id_router_028_src_endofpacket;                                                           // id_router_028:src_endofpacket -> width_adapter_045:in_endofpacket
	wire         id_router_028_src_valid;                                                                 // id_router_028:src_valid -> width_adapter_045:in_valid
	wire         id_router_028_src_startofpacket;                                                         // id_router_028:src_startofpacket -> width_adapter_045:in_startofpacket
	wire  [65:0] id_router_028_src_data;                                                                  // id_router_028:src_data -> width_adapter_045:in_data
	wire  [57:0] id_router_028_src_channel;                                                               // id_router_028:src_channel -> width_adapter_045:in_channel
	wire         id_router_028_src_ready;                                                                 // width_adapter_045:in_ready -> id_router_028:src_ready
	wire         width_adapter_045_src_endofpacket;                                                       // width_adapter_045:out_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	wire         width_adapter_045_src_valid;                                                             // width_adapter_045:out_valid -> rsp_xbar_demux_028:sink_valid
	wire         width_adapter_045_src_startofpacket;                                                     // width_adapter_045:out_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	wire  [92:0] width_adapter_045_src_data;                                                              // width_adapter_045:out_data -> rsp_xbar_demux_028:sink_data
	wire         width_adapter_045_src_ready;                                                             // rsp_xbar_demux_028:sink_ready -> width_adapter_045:out_ready
	wire  [57:0] width_adapter_045_src_channel;                                                           // width_adapter_045:out_channel -> rsp_xbar_demux_028:sink_channel
	wire         cmd_xbar_demux_src29_ready;                                                              // width_adapter_046:in_ready -> cmd_xbar_demux:src29_ready
	wire         width_adapter_046_src_endofpacket;                                                       // width_adapter_046:out_endofpacket -> burst_adapter_050:sink0_endofpacket
	wire         width_adapter_046_src_valid;                                                             // width_adapter_046:out_valid -> burst_adapter_050:sink0_valid
	wire         width_adapter_046_src_startofpacket;                                                     // width_adapter_046:out_startofpacket -> burst_adapter_050:sink0_startofpacket
	wire  [65:0] width_adapter_046_src_data;                                                              // width_adapter_046:out_data -> burst_adapter_050:sink0_data
	wire         width_adapter_046_src_ready;                                                             // burst_adapter_050:sink0_ready -> width_adapter_046:out_ready
	wire  [57:0] width_adapter_046_src_channel;                                                           // width_adapter_046:out_channel -> burst_adapter_050:sink0_channel
	wire         id_router_029_src_endofpacket;                                                           // id_router_029:src_endofpacket -> width_adapter_047:in_endofpacket
	wire         id_router_029_src_valid;                                                                 // id_router_029:src_valid -> width_adapter_047:in_valid
	wire         id_router_029_src_startofpacket;                                                         // id_router_029:src_startofpacket -> width_adapter_047:in_startofpacket
	wire  [65:0] id_router_029_src_data;                                                                  // id_router_029:src_data -> width_adapter_047:in_data
	wire  [57:0] id_router_029_src_channel;                                                               // id_router_029:src_channel -> width_adapter_047:in_channel
	wire         id_router_029_src_ready;                                                                 // width_adapter_047:in_ready -> id_router_029:src_ready
	wire         width_adapter_047_src_endofpacket;                                                       // width_adapter_047:out_endofpacket -> rsp_xbar_demux_029:sink_endofpacket
	wire         width_adapter_047_src_valid;                                                             // width_adapter_047:out_valid -> rsp_xbar_demux_029:sink_valid
	wire         width_adapter_047_src_startofpacket;                                                     // width_adapter_047:out_startofpacket -> rsp_xbar_demux_029:sink_startofpacket
	wire  [92:0] width_adapter_047_src_data;                                                              // width_adapter_047:out_data -> rsp_xbar_demux_029:sink_data
	wire         width_adapter_047_src_ready;                                                             // rsp_xbar_demux_029:sink_ready -> width_adapter_047:out_ready
	wire  [57:0] width_adapter_047_src_channel;                                                           // width_adapter_047:out_channel -> rsp_xbar_demux_029:sink_channel
	wire         cmd_xbar_demux_src30_ready;                                                              // width_adapter_048:in_ready -> cmd_xbar_demux:src30_ready
	wire         width_adapter_048_src_endofpacket;                                                       // width_adapter_048:out_endofpacket -> burst_adapter_019:sink0_endofpacket
	wire         width_adapter_048_src_valid;                                                             // width_adapter_048:out_valid -> burst_adapter_019:sink0_valid
	wire         width_adapter_048_src_startofpacket;                                                     // width_adapter_048:out_startofpacket -> burst_adapter_019:sink0_startofpacket
	wire  [65:0] width_adapter_048_src_data;                                                              // width_adapter_048:out_data -> burst_adapter_019:sink0_data
	wire         width_adapter_048_src_ready;                                                             // burst_adapter_019:sink0_ready -> width_adapter_048:out_ready
	wire  [57:0] width_adapter_048_src_channel;                                                           // width_adapter_048:out_channel -> burst_adapter_019:sink0_channel
	wire         id_router_030_src_endofpacket;                                                           // id_router_030:src_endofpacket -> width_adapter_049:in_endofpacket
	wire         id_router_030_src_valid;                                                                 // id_router_030:src_valid -> width_adapter_049:in_valid
	wire         id_router_030_src_startofpacket;                                                         // id_router_030:src_startofpacket -> width_adapter_049:in_startofpacket
	wire  [65:0] id_router_030_src_data;                                                                  // id_router_030:src_data -> width_adapter_049:in_data
	wire  [57:0] id_router_030_src_channel;                                                               // id_router_030:src_channel -> width_adapter_049:in_channel
	wire         id_router_030_src_ready;                                                                 // width_adapter_049:in_ready -> id_router_030:src_ready
	wire         width_adapter_049_src_endofpacket;                                                       // width_adapter_049:out_endofpacket -> rsp_xbar_demux_030:sink_endofpacket
	wire         width_adapter_049_src_valid;                                                             // width_adapter_049:out_valid -> rsp_xbar_demux_030:sink_valid
	wire         width_adapter_049_src_startofpacket;                                                     // width_adapter_049:out_startofpacket -> rsp_xbar_demux_030:sink_startofpacket
	wire  [92:0] width_adapter_049_src_data;                                                              // width_adapter_049:out_data -> rsp_xbar_demux_030:sink_data
	wire         width_adapter_049_src_ready;                                                             // rsp_xbar_demux_030:sink_ready -> width_adapter_049:out_ready
	wire  [57:0] width_adapter_049_src_channel;                                                           // width_adapter_049:out_channel -> rsp_xbar_demux_030:sink_channel
	wire         cmd_xbar_demux_src31_ready;                                                              // width_adapter_050:in_ready -> cmd_xbar_demux:src31_ready
	wire         width_adapter_050_src_endofpacket;                                                       // width_adapter_050:out_endofpacket -> burst_adapter_021:sink0_endofpacket
	wire         width_adapter_050_src_valid;                                                             // width_adapter_050:out_valid -> burst_adapter_021:sink0_valid
	wire         width_adapter_050_src_startofpacket;                                                     // width_adapter_050:out_startofpacket -> burst_adapter_021:sink0_startofpacket
	wire  [65:0] width_adapter_050_src_data;                                                              // width_adapter_050:out_data -> burst_adapter_021:sink0_data
	wire         width_adapter_050_src_ready;                                                             // burst_adapter_021:sink0_ready -> width_adapter_050:out_ready
	wire  [57:0] width_adapter_050_src_channel;                                                           // width_adapter_050:out_channel -> burst_adapter_021:sink0_channel
	wire         id_router_031_src_endofpacket;                                                           // id_router_031:src_endofpacket -> width_adapter_051:in_endofpacket
	wire         id_router_031_src_valid;                                                                 // id_router_031:src_valid -> width_adapter_051:in_valid
	wire         id_router_031_src_startofpacket;                                                         // id_router_031:src_startofpacket -> width_adapter_051:in_startofpacket
	wire  [65:0] id_router_031_src_data;                                                                  // id_router_031:src_data -> width_adapter_051:in_data
	wire  [57:0] id_router_031_src_channel;                                                               // id_router_031:src_channel -> width_adapter_051:in_channel
	wire         id_router_031_src_ready;                                                                 // width_adapter_051:in_ready -> id_router_031:src_ready
	wire         width_adapter_051_src_endofpacket;                                                       // width_adapter_051:out_endofpacket -> rsp_xbar_demux_031:sink_endofpacket
	wire         width_adapter_051_src_valid;                                                             // width_adapter_051:out_valid -> rsp_xbar_demux_031:sink_valid
	wire         width_adapter_051_src_startofpacket;                                                     // width_adapter_051:out_startofpacket -> rsp_xbar_demux_031:sink_startofpacket
	wire  [92:0] width_adapter_051_src_data;                                                              // width_adapter_051:out_data -> rsp_xbar_demux_031:sink_data
	wire         width_adapter_051_src_ready;                                                             // rsp_xbar_demux_031:sink_ready -> width_adapter_051:out_ready
	wire  [57:0] width_adapter_051_src_channel;                                                           // width_adapter_051:out_channel -> rsp_xbar_demux_031:sink_channel
	wire         cmd_xbar_demux_src32_ready;                                                              // width_adapter_052:in_ready -> cmd_xbar_demux:src32_ready
	wire         width_adapter_052_src_endofpacket;                                                       // width_adapter_052:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire         width_adapter_052_src_valid;                                                             // width_adapter_052:out_valid -> burst_adapter:sink0_valid
	wire         width_adapter_052_src_startofpacket;                                                     // width_adapter_052:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [65:0] width_adapter_052_src_data;                                                              // width_adapter_052:out_data -> burst_adapter:sink0_data
	wire         width_adapter_052_src_ready;                                                             // burst_adapter:sink0_ready -> width_adapter_052:out_ready
	wire  [57:0] width_adapter_052_src_channel;                                                           // width_adapter_052:out_channel -> burst_adapter:sink0_channel
	wire         id_router_032_src_endofpacket;                                                           // id_router_032:src_endofpacket -> width_adapter_053:in_endofpacket
	wire         id_router_032_src_valid;                                                                 // id_router_032:src_valid -> width_adapter_053:in_valid
	wire         id_router_032_src_startofpacket;                                                         // id_router_032:src_startofpacket -> width_adapter_053:in_startofpacket
	wire  [65:0] id_router_032_src_data;                                                                  // id_router_032:src_data -> width_adapter_053:in_data
	wire  [57:0] id_router_032_src_channel;                                                               // id_router_032:src_channel -> width_adapter_053:in_channel
	wire         id_router_032_src_ready;                                                                 // width_adapter_053:in_ready -> id_router_032:src_ready
	wire         width_adapter_053_src_endofpacket;                                                       // width_adapter_053:out_endofpacket -> rsp_xbar_demux_032:sink_endofpacket
	wire         width_adapter_053_src_valid;                                                             // width_adapter_053:out_valid -> rsp_xbar_demux_032:sink_valid
	wire         width_adapter_053_src_startofpacket;                                                     // width_adapter_053:out_startofpacket -> rsp_xbar_demux_032:sink_startofpacket
	wire  [92:0] width_adapter_053_src_data;                                                              // width_adapter_053:out_data -> rsp_xbar_demux_032:sink_data
	wire         width_adapter_053_src_ready;                                                             // rsp_xbar_demux_032:sink_ready -> width_adapter_053:out_ready
	wire  [57:0] width_adapter_053_src_channel;                                                           // width_adapter_053:out_channel -> rsp_xbar_demux_032:sink_channel
	wire         cmd_xbar_demux_src33_ready;                                                              // width_adapter_054:in_ready -> cmd_xbar_demux:src33_ready
	wire         width_adapter_054_src_endofpacket;                                                       // width_adapter_054:out_endofpacket -> burst_adapter_009:sink0_endofpacket
	wire         width_adapter_054_src_valid;                                                             // width_adapter_054:out_valid -> burst_adapter_009:sink0_valid
	wire         width_adapter_054_src_startofpacket;                                                     // width_adapter_054:out_startofpacket -> burst_adapter_009:sink0_startofpacket
	wire  [65:0] width_adapter_054_src_data;                                                              // width_adapter_054:out_data -> burst_adapter_009:sink0_data
	wire         width_adapter_054_src_ready;                                                             // burst_adapter_009:sink0_ready -> width_adapter_054:out_ready
	wire  [57:0] width_adapter_054_src_channel;                                                           // width_adapter_054:out_channel -> burst_adapter_009:sink0_channel
	wire         id_router_033_src_endofpacket;                                                           // id_router_033:src_endofpacket -> width_adapter_055:in_endofpacket
	wire         id_router_033_src_valid;                                                                 // id_router_033:src_valid -> width_adapter_055:in_valid
	wire         id_router_033_src_startofpacket;                                                         // id_router_033:src_startofpacket -> width_adapter_055:in_startofpacket
	wire  [65:0] id_router_033_src_data;                                                                  // id_router_033:src_data -> width_adapter_055:in_data
	wire  [57:0] id_router_033_src_channel;                                                               // id_router_033:src_channel -> width_adapter_055:in_channel
	wire         id_router_033_src_ready;                                                                 // width_adapter_055:in_ready -> id_router_033:src_ready
	wire         width_adapter_055_src_endofpacket;                                                       // width_adapter_055:out_endofpacket -> rsp_xbar_demux_033:sink_endofpacket
	wire         width_adapter_055_src_valid;                                                             // width_adapter_055:out_valid -> rsp_xbar_demux_033:sink_valid
	wire         width_adapter_055_src_startofpacket;                                                     // width_adapter_055:out_startofpacket -> rsp_xbar_demux_033:sink_startofpacket
	wire  [92:0] width_adapter_055_src_data;                                                              // width_adapter_055:out_data -> rsp_xbar_demux_033:sink_data
	wire         width_adapter_055_src_ready;                                                             // rsp_xbar_demux_033:sink_ready -> width_adapter_055:out_ready
	wire  [57:0] width_adapter_055_src_channel;                                                           // width_adapter_055:out_channel -> rsp_xbar_demux_033:sink_channel
	wire         cmd_xbar_demux_src34_ready;                                                              // width_adapter_056:in_ready -> cmd_xbar_demux:src34_ready
	wire         width_adapter_056_src_endofpacket;                                                       // width_adapter_056:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire         width_adapter_056_src_valid;                                                             // width_adapter_056:out_valid -> burst_adapter_001:sink0_valid
	wire         width_adapter_056_src_startofpacket;                                                     // width_adapter_056:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [65:0] width_adapter_056_src_data;                                                              // width_adapter_056:out_data -> burst_adapter_001:sink0_data
	wire         width_adapter_056_src_ready;                                                             // burst_adapter_001:sink0_ready -> width_adapter_056:out_ready
	wire  [57:0] width_adapter_056_src_channel;                                                           // width_adapter_056:out_channel -> burst_adapter_001:sink0_channel
	wire         id_router_034_src_endofpacket;                                                           // id_router_034:src_endofpacket -> width_adapter_057:in_endofpacket
	wire         id_router_034_src_valid;                                                                 // id_router_034:src_valid -> width_adapter_057:in_valid
	wire         id_router_034_src_startofpacket;                                                         // id_router_034:src_startofpacket -> width_adapter_057:in_startofpacket
	wire  [65:0] id_router_034_src_data;                                                                  // id_router_034:src_data -> width_adapter_057:in_data
	wire  [57:0] id_router_034_src_channel;                                                               // id_router_034:src_channel -> width_adapter_057:in_channel
	wire         id_router_034_src_ready;                                                                 // width_adapter_057:in_ready -> id_router_034:src_ready
	wire         width_adapter_057_src_endofpacket;                                                       // width_adapter_057:out_endofpacket -> rsp_xbar_demux_034:sink_endofpacket
	wire         width_adapter_057_src_valid;                                                             // width_adapter_057:out_valid -> rsp_xbar_demux_034:sink_valid
	wire         width_adapter_057_src_startofpacket;                                                     // width_adapter_057:out_startofpacket -> rsp_xbar_demux_034:sink_startofpacket
	wire  [92:0] width_adapter_057_src_data;                                                              // width_adapter_057:out_data -> rsp_xbar_demux_034:sink_data
	wire         width_adapter_057_src_ready;                                                             // rsp_xbar_demux_034:sink_ready -> width_adapter_057:out_ready
	wire  [57:0] width_adapter_057_src_channel;                                                           // width_adapter_057:out_channel -> rsp_xbar_demux_034:sink_channel
	wire         cmd_xbar_demux_src35_ready;                                                              // width_adapter_058:in_ready -> cmd_xbar_demux:src35_ready
	wire         width_adapter_058_src_endofpacket;                                                       // width_adapter_058:out_endofpacket -> burst_adapter_044:sink0_endofpacket
	wire         width_adapter_058_src_valid;                                                             // width_adapter_058:out_valid -> burst_adapter_044:sink0_valid
	wire         width_adapter_058_src_startofpacket;                                                     // width_adapter_058:out_startofpacket -> burst_adapter_044:sink0_startofpacket
	wire  [65:0] width_adapter_058_src_data;                                                              // width_adapter_058:out_data -> burst_adapter_044:sink0_data
	wire         width_adapter_058_src_ready;                                                             // burst_adapter_044:sink0_ready -> width_adapter_058:out_ready
	wire  [57:0] width_adapter_058_src_channel;                                                           // width_adapter_058:out_channel -> burst_adapter_044:sink0_channel
	wire         id_router_035_src_endofpacket;                                                           // id_router_035:src_endofpacket -> width_adapter_059:in_endofpacket
	wire         id_router_035_src_valid;                                                                 // id_router_035:src_valid -> width_adapter_059:in_valid
	wire         id_router_035_src_startofpacket;                                                         // id_router_035:src_startofpacket -> width_adapter_059:in_startofpacket
	wire  [65:0] id_router_035_src_data;                                                                  // id_router_035:src_data -> width_adapter_059:in_data
	wire  [57:0] id_router_035_src_channel;                                                               // id_router_035:src_channel -> width_adapter_059:in_channel
	wire         id_router_035_src_ready;                                                                 // width_adapter_059:in_ready -> id_router_035:src_ready
	wire         width_adapter_059_src_endofpacket;                                                       // width_adapter_059:out_endofpacket -> rsp_xbar_demux_035:sink_endofpacket
	wire         width_adapter_059_src_valid;                                                             // width_adapter_059:out_valid -> rsp_xbar_demux_035:sink_valid
	wire         width_adapter_059_src_startofpacket;                                                     // width_adapter_059:out_startofpacket -> rsp_xbar_demux_035:sink_startofpacket
	wire  [92:0] width_adapter_059_src_data;                                                              // width_adapter_059:out_data -> rsp_xbar_demux_035:sink_data
	wire         width_adapter_059_src_ready;                                                             // rsp_xbar_demux_035:sink_ready -> width_adapter_059:out_ready
	wire  [57:0] width_adapter_059_src_channel;                                                           // width_adapter_059:out_channel -> rsp_xbar_demux_035:sink_channel
	wire         cmd_xbar_demux_src36_ready;                                                              // width_adapter_060:in_ready -> cmd_xbar_demux:src36_ready
	wire         width_adapter_060_src_endofpacket;                                                       // width_adapter_060:out_endofpacket -> burst_adapter_041:sink0_endofpacket
	wire         width_adapter_060_src_valid;                                                             // width_adapter_060:out_valid -> burst_adapter_041:sink0_valid
	wire         width_adapter_060_src_startofpacket;                                                     // width_adapter_060:out_startofpacket -> burst_adapter_041:sink0_startofpacket
	wire  [65:0] width_adapter_060_src_data;                                                              // width_adapter_060:out_data -> burst_adapter_041:sink0_data
	wire         width_adapter_060_src_ready;                                                             // burst_adapter_041:sink0_ready -> width_adapter_060:out_ready
	wire  [57:0] width_adapter_060_src_channel;                                                           // width_adapter_060:out_channel -> burst_adapter_041:sink0_channel
	wire         id_router_036_src_endofpacket;                                                           // id_router_036:src_endofpacket -> width_adapter_061:in_endofpacket
	wire         id_router_036_src_valid;                                                                 // id_router_036:src_valid -> width_adapter_061:in_valid
	wire         id_router_036_src_startofpacket;                                                         // id_router_036:src_startofpacket -> width_adapter_061:in_startofpacket
	wire  [65:0] id_router_036_src_data;                                                                  // id_router_036:src_data -> width_adapter_061:in_data
	wire  [57:0] id_router_036_src_channel;                                                               // id_router_036:src_channel -> width_adapter_061:in_channel
	wire         id_router_036_src_ready;                                                                 // width_adapter_061:in_ready -> id_router_036:src_ready
	wire         width_adapter_061_src_endofpacket;                                                       // width_adapter_061:out_endofpacket -> rsp_xbar_demux_036:sink_endofpacket
	wire         width_adapter_061_src_valid;                                                             // width_adapter_061:out_valid -> rsp_xbar_demux_036:sink_valid
	wire         width_adapter_061_src_startofpacket;                                                     // width_adapter_061:out_startofpacket -> rsp_xbar_demux_036:sink_startofpacket
	wire  [92:0] width_adapter_061_src_data;                                                              // width_adapter_061:out_data -> rsp_xbar_demux_036:sink_data
	wire         width_adapter_061_src_ready;                                                             // rsp_xbar_demux_036:sink_ready -> width_adapter_061:out_ready
	wire  [57:0] width_adapter_061_src_channel;                                                           // width_adapter_061:out_channel -> rsp_xbar_demux_036:sink_channel
	wire         cmd_xbar_demux_src37_ready;                                                              // width_adapter_062:in_ready -> cmd_xbar_demux:src37_ready
	wire         width_adapter_062_src_endofpacket;                                                       // width_adapter_062:out_endofpacket -> burst_adapter_031:sink0_endofpacket
	wire         width_adapter_062_src_valid;                                                             // width_adapter_062:out_valid -> burst_adapter_031:sink0_valid
	wire         width_adapter_062_src_startofpacket;                                                     // width_adapter_062:out_startofpacket -> burst_adapter_031:sink0_startofpacket
	wire  [65:0] width_adapter_062_src_data;                                                              // width_adapter_062:out_data -> burst_adapter_031:sink0_data
	wire         width_adapter_062_src_ready;                                                             // burst_adapter_031:sink0_ready -> width_adapter_062:out_ready
	wire  [57:0] width_adapter_062_src_channel;                                                           // width_adapter_062:out_channel -> burst_adapter_031:sink0_channel
	wire         id_router_037_src_endofpacket;                                                           // id_router_037:src_endofpacket -> width_adapter_063:in_endofpacket
	wire         id_router_037_src_valid;                                                                 // id_router_037:src_valid -> width_adapter_063:in_valid
	wire         id_router_037_src_startofpacket;                                                         // id_router_037:src_startofpacket -> width_adapter_063:in_startofpacket
	wire  [65:0] id_router_037_src_data;                                                                  // id_router_037:src_data -> width_adapter_063:in_data
	wire  [57:0] id_router_037_src_channel;                                                               // id_router_037:src_channel -> width_adapter_063:in_channel
	wire         id_router_037_src_ready;                                                                 // width_adapter_063:in_ready -> id_router_037:src_ready
	wire         width_adapter_063_src_endofpacket;                                                       // width_adapter_063:out_endofpacket -> rsp_xbar_demux_037:sink_endofpacket
	wire         width_adapter_063_src_valid;                                                             // width_adapter_063:out_valid -> rsp_xbar_demux_037:sink_valid
	wire         width_adapter_063_src_startofpacket;                                                     // width_adapter_063:out_startofpacket -> rsp_xbar_demux_037:sink_startofpacket
	wire  [92:0] width_adapter_063_src_data;                                                              // width_adapter_063:out_data -> rsp_xbar_demux_037:sink_data
	wire         width_adapter_063_src_ready;                                                             // rsp_xbar_demux_037:sink_ready -> width_adapter_063:out_ready
	wire  [57:0] width_adapter_063_src_channel;                                                           // width_adapter_063:out_channel -> rsp_xbar_demux_037:sink_channel
	wire         cmd_xbar_demux_src38_ready;                                                              // width_adapter_064:in_ready -> cmd_xbar_demux:src38_ready
	wire         width_adapter_064_src_endofpacket;                                                       // width_adapter_064:out_endofpacket -> burst_adapter_026:sink0_endofpacket
	wire         width_adapter_064_src_valid;                                                             // width_adapter_064:out_valid -> burst_adapter_026:sink0_valid
	wire         width_adapter_064_src_startofpacket;                                                     // width_adapter_064:out_startofpacket -> burst_adapter_026:sink0_startofpacket
	wire  [65:0] width_adapter_064_src_data;                                                              // width_adapter_064:out_data -> burst_adapter_026:sink0_data
	wire         width_adapter_064_src_ready;                                                             // burst_adapter_026:sink0_ready -> width_adapter_064:out_ready
	wire  [57:0] width_adapter_064_src_channel;                                                           // width_adapter_064:out_channel -> burst_adapter_026:sink0_channel
	wire         id_router_038_src_endofpacket;                                                           // id_router_038:src_endofpacket -> width_adapter_065:in_endofpacket
	wire         id_router_038_src_valid;                                                                 // id_router_038:src_valid -> width_adapter_065:in_valid
	wire         id_router_038_src_startofpacket;                                                         // id_router_038:src_startofpacket -> width_adapter_065:in_startofpacket
	wire  [65:0] id_router_038_src_data;                                                                  // id_router_038:src_data -> width_adapter_065:in_data
	wire  [57:0] id_router_038_src_channel;                                                               // id_router_038:src_channel -> width_adapter_065:in_channel
	wire         id_router_038_src_ready;                                                                 // width_adapter_065:in_ready -> id_router_038:src_ready
	wire         width_adapter_065_src_endofpacket;                                                       // width_adapter_065:out_endofpacket -> rsp_xbar_demux_038:sink_endofpacket
	wire         width_adapter_065_src_valid;                                                             // width_adapter_065:out_valid -> rsp_xbar_demux_038:sink_valid
	wire         width_adapter_065_src_startofpacket;                                                     // width_adapter_065:out_startofpacket -> rsp_xbar_demux_038:sink_startofpacket
	wire  [92:0] width_adapter_065_src_data;                                                              // width_adapter_065:out_data -> rsp_xbar_demux_038:sink_data
	wire         width_adapter_065_src_ready;                                                             // rsp_xbar_demux_038:sink_ready -> width_adapter_065:out_ready
	wire  [57:0] width_adapter_065_src_channel;                                                           // width_adapter_065:out_channel -> rsp_xbar_demux_038:sink_channel
	wire         cmd_xbar_demux_src39_ready;                                                              // width_adapter_066:in_ready -> cmd_xbar_demux:src39_ready
	wire         width_adapter_066_src_endofpacket;                                                       // width_adapter_066:out_endofpacket -> burst_adapter_017:sink0_endofpacket
	wire         width_adapter_066_src_valid;                                                             // width_adapter_066:out_valid -> burst_adapter_017:sink0_valid
	wire         width_adapter_066_src_startofpacket;                                                     // width_adapter_066:out_startofpacket -> burst_adapter_017:sink0_startofpacket
	wire  [65:0] width_adapter_066_src_data;                                                              // width_adapter_066:out_data -> burst_adapter_017:sink0_data
	wire         width_adapter_066_src_ready;                                                             // burst_adapter_017:sink0_ready -> width_adapter_066:out_ready
	wire  [57:0] width_adapter_066_src_channel;                                                           // width_adapter_066:out_channel -> burst_adapter_017:sink0_channel
	wire         id_router_039_src_endofpacket;                                                           // id_router_039:src_endofpacket -> width_adapter_067:in_endofpacket
	wire         id_router_039_src_valid;                                                                 // id_router_039:src_valid -> width_adapter_067:in_valid
	wire         id_router_039_src_startofpacket;                                                         // id_router_039:src_startofpacket -> width_adapter_067:in_startofpacket
	wire  [65:0] id_router_039_src_data;                                                                  // id_router_039:src_data -> width_adapter_067:in_data
	wire  [57:0] id_router_039_src_channel;                                                               // id_router_039:src_channel -> width_adapter_067:in_channel
	wire         id_router_039_src_ready;                                                                 // width_adapter_067:in_ready -> id_router_039:src_ready
	wire         width_adapter_067_src_endofpacket;                                                       // width_adapter_067:out_endofpacket -> rsp_xbar_demux_039:sink_endofpacket
	wire         width_adapter_067_src_valid;                                                             // width_adapter_067:out_valid -> rsp_xbar_demux_039:sink_valid
	wire         width_adapter_067_src_startofpacket;                                                     // width_adapter_067:out_startofpacket -> rsp_xbar_demux_039:sink_startofpacket
	wire  [92:0] width_adapter_067_src_data;                                                              // width_adapter_067:out_data -> rsp_xbar_demux_039:sink_data
	wire         width_adapter_067_src_ready;                                                             // rsp_xbar_demux_039:sink_ready -> width_adapter_067:out_ready
	wire  [57:0] width_adapter_067_src_channel;                                                           // width_adapter_067:out_channel -> rsp_xbar_demux_039:sink_channel
	wire         cmd_xbar_demux_src40_ready;                                                              // width_adapter_068:in_ready -> cmd_xbar_demux:src40_ready
	wire         width_adapter_068_src_endofpacket;                                                       // width_adapter_068:out_endofpacket -> burst_adapter_015:sink0_endofpacket
	wire         width_adapter_068_src_valid;                                                             // width_adapter_068:out_valid -> burst_adapter_015:sink0_valid
	wire         width_adapter_068_src_startofpacket;                                                     // width_adapter_068:out_startofpacket -> burst_adapter_015:sink0_startofpacket
	wire  [65:0] width_adapter_068_src_data;                                                              // width_adapter_068:out_data -> burst_adapter_015:sink0_data
	wire         width_adapter_068_src_ready;                                                             // burst_adapter_015:sink0_ready -> width_adapter_068:out_ready
	wire  [57:0] width_adapter_068_src_channel;                                                           // width_adapter_068:out_channel -> burst_adapter_015:sink0_channel
	wire         id_router_040_src_endofpacket;                                                           // id_router_040:src_endofpacket -> width_adapter_069:in_endofpacket
	wire         id_router_040_src_valid;                                                                 // id_router_040:src_valid -> width_adapter_069:in_valid
	wire         id_router_040_src_startofpacket;                                                         // id_router_040:src_startofpacket -> width_adapter_069:in_startofpacket
	wire  [65:0] id_router_040_src_data;                                                                  // id_router_040:src_data -> width_adapter_069:in_data
	wire  [57:0] id_router_040_src_channel;                                                               // id_router_040:src_channel -> width_adapter_069:in_channel
	wire         id_router_040_src_ready;                                                                 // width_adapter_069:in_ready -> id_router_040:src_ready
	wire         width_adapter_069_src_endofpacket;                                                       // width_adapter_069:out_endofpacket -> rsp_xbar_demux_040:sink_endofpacket
	wire         width_adapter_069_src_valid;                                                             // width_adapter_069:out_valid -> rsp_xbar_demux_040:sink_valid
	wire         width_adapter_069_src_startofpacket;                                                     // width_adapter_069:out_startofpacket -> rsp_xbar_demux_040:sink_startofpacket
	wire  [92:0] width_adapter_069_src_data;                                                              // width_adapter_069:out_data -> rsp_xbar_demux_040:sink_data
	wire         width_adapter_069_src_ready;                                                             // rsp_xbar_demux_040:sink_ready -> width_adapter_069:out_ready
	wire  [57:0] width_adapter_069_src_channel;                                                           // width_adapter_069:out_channel -> rsp_xbar_demux_040:sink_channel
	wire         cmd_xbar_demux_src41_ready;                                                              // width_adapter_070:in_ready -> cmd_xbar_demux:src41_ready
	wire         width_adapter_070_src_endofpacket;                                                       // width_adapter_070:out_endofpacket -> burst_adapter_032:sink0_endofpacket
	wire         width_adapter_070_src_valid;                                                             // width_adapter_070:out_valid -> burst_adapter_032:sink0_valid
	wire         width_adapter_070_src_startofpacket;                                                     // width_adapter_070:out_startofpacket -> burst_adapter_032:sink0_startofpacket
	wire  [65:0] width_adapter_070_src_data;                                                              // width_adapter_070:out_data -> burst_adapter_032:sink0_data
	wire         width_adapter_070_src_ready;                                                             // burst_adapter_032:sink0_ready -> width_adapter_070:out_ready
	wire  [57:0] width_adapter_070_src_channel;                                                           // width_adapter_070:out_channel -> burst_adapter_032:sink0_channel
	wire         id_router_041_src_endofpacket;                                                           // id_router_041:src_endofpacket -> width_adapter_071:in_endofpacket
	wire         id_router_041_src_valid;                                                                 // id_router_041:src_valid -> width_adapter_071:in_valid
	wire         id_router_041_src_startofpacket;                                                         // id_router_041:src_startofpacket -> width_adapter_071:in_startofpacket
	wire  [65:0] id_router_041_src_data;                                                                  // id_router_041:src_data -> width_adapter_071:in_data
	wire  [57:0] id_router_041_src_channel;                                                               // id_router_041:src_channel -> width_adapter_071:in_channel
	wire         id_router_041_src_ready;                                                                 // width_adapter_071:in_ready -> id_router_041:src_ready
	wire         width_adapter_071_src_endofpacket;                                                       // width_adapter_071:out_endofpacket -> rsp_xbar_demux_041:sink_endofpacket
	wire         width_adapter_071_src_valid;                                                             // width_adapter_071:out_valid -> rsp_xbar_demux_041:sink_valid
	wire         width_adapter_071_src_startofpacket;                                                     // width_adapter_071:out_startofpacket -> rsp_xbar_demux_041:sink_startofpacket
	wire  [92:0] width_adapter_071_src_data;                                                              // width_adapter_071:out_data -> rsp_xbar_demux_041:sink_data
	wire         width_adapter_071_src_ready;                                                             // rsp_xbar_demux_041:sink_ready -> width_adapter_071:out_ready
	wire  [57:0] width_adapter_071_src_channel;                                                           // width_adapter_071:out_channel -> rsp_xbar_demux_041:sink_channel
	wire         cmd_xbar_demux_src42_ready;                                                              // width_adapter_072:in_ready -> cmd_xbar_demux:src42_ready
	wire         width_adapter_072_src_endofpacket;                                                       // width_adapter_072:out_endofpacket -> burst_adapter_028:sink0_endofpacket
	wire         width_adapter_072_src_valid;                                                             // width_adapter_072:out_valid -> burst_adapter_028:sink0_valid
	wire         width_adapter_072_src_startofpacket;                                                     // width_adapter_072:out_startofpacket -> burst_adapter_028:sink0_startofpacket
	wire  [65:0] width_adapter_072_src_data;                                                              // width_adapter_072:out_data -> burst_adapter_028:sink0_data
	wire         width_adapter_072_src_ready;                                                             // burst_adapter_028:sink0_ready -> width_adapter_072:out_ready
	wire  [57:0] width_adapter_072_src_channel;                                                           // width_adapter_072:out_channel -> burst_adapter_028:sink0_channel
	wire         id_router_042_src_endofpacket;                                                           // id_router_042:src_endofpacket -> width_adapter_073:in_endofpacket
	wire         id_router_042_src_valid;                                                                 // id_router_042:src_valid -> width_adapter_073:in_valid
	wire         id_router_042_src_startofpacket;                                                         // id_router_042:src_startofpacket -> width_adapter_073:in_startofpacket
	wire  [65:0] id_router_042_src_data;                                                                  // id_router_042:src_data -> width_adapter_073:in_data
	wire  [57:0] id_router_042_src_channel;                                                               // id_router_042:src_channel -> width_adapter_073:in_channel
	wire         id_router_042_src_ready;                                                                 // width_adapter_073:in_ready -> id_router_042:src_ready
	wire         width_adapter_073_src_endofpacket;                                                       // width_adapter_073:out_endofpacket -> rsp_xbar_demux_042:sink_endofpacket
	wire         width_adapter_073_src_valid;                                                             // width_adapter_073:out_valid -> rsp_xbar_demux_042:sink_valid
	wire         width_adapter_073_src_startofpacket;                                                     // width_adapter_073:out_startofpacket -> rsp_xbar_demux_042:sink_startofpacket
	wire  [92:0] width_adapter_073_src_data;                                                              // width_adapter_073:out_data -> rsp_xbar_demux_042:sink_data
	wire         width_adapter_073_src_ready;                                                             // rsp_xbar_demux_042:sink_ready -> width_adapter_073:out_ready
	wire  [57:0] width_adapter_073_src_channel;                                                           // width_adapter_073:out_channel -> rsp_xbar_demux_042:sink_channel
	wire         cmd_xbar_demux_src43_ready;                                                              // width_adapter_074:in_ready -> cmd_xbar_demux:src43_ready
	wire         width_adapter_074_src_endofpacket;                                                       // width_adapter_074:out_endofpacket -> burst_adapter_013:sink0_endofpacket
	wire         width_adapter_074_src_valid;                                                             // width_adapter_074:out_valid -> burst_adapter_013:sink0_valid
	wire         width_adapter_074_src_startofpacket;                                                     // width_adapter_074:out_startofpacket -> burst_adapter_013:sink0_startofpacket
	wire  [65:0] width_adapter_074_src_data;                                                              // width_adapter_074:out_data -> burst_adapter_013:sink0_data
	wire         width_adapter_074_src_ready;                                                             // burst_adapter_013:sink0_ready -> width_adapter_074:out_ready
	wire  [57:0] width_adapter_074_src_channel;                                                           // width_adapter_074:out_channel -> burst_adapter_013:sink0_channel
	wire         id_router_043_src_endofpacket;                                                           // id_router_043:src_endofpacket -> width_adapter_075:in_endofpacket
	wire         id_router_043_src_valid;                                                                 // id_router_043:src_valid -> width_adapter_075:in_valid
	wire         id_router_043_src_startofpacket;                                                         // id_router_043:src_startofpacket -> width_adapter_075:in_startofpacket
	wire  [65:0] id_router_043_src_data;                                                                  // id_router_043:src_data -> width_adapter_075:in_data
	wire  [57:0] id_router_043_src_channel;                                                               // id_router_043:src_channel -> width_adapter_075:in_channel
	wire         id_router_043_src_ready;                                                                 // width_adapter_075:in_ready -> id_router_043:src_ready
	wire         width_adapter_075_src_endofpacket;                                                       // width_adapter_075:out_endofpacket -> rsp_xbar_demux_043:sink_endofpacket
	wire         width_adapter_075_src_valid;                                                             // width_adapter_075:out_valid -> rsp_xbar_demux_043:sink_valid
	wire         width_adapter_075_src_startofpacket;                                                     // width_adapter_075:out_startofpacket -> rsp_xbar_demux_043:sink_startofpacket
	wire  [92:0] width_adapter_075_src_data;                                                              // width_adapter_075:out_data -> rsp_xbar_demux_043:sink_data
	wire         width_adapter_075_src_ready;                                                             // rsp_xbar_demux_043:sink_ready -> width_adapter_075:out_ready
	wire  [57:0] width_adapter_075_src_channel;                                                           // width_adapter_075:out_channel -> rsp_xbar_demux_043:sink_channel
	wire         cmd_xbar_demux_src44_ready;                                                              // width_adapter_076:in_ready -> cmd_xbar_demux:src44_ready
	wire         width_adapter_076_src_endofpacket;                                                       // width_adapter_076:out_endofpacket -> burst_adapter_029:sink0_endofpacket
	wire         width_adapter_076_src_valid;                                                             // width_adapter_076:out_valid -> burst_adapter_029:sink0_valid
	wire         width_adapter_076_src_startofpacket;                                                     // width_adapter_076:out_startofpacket -> burst_adapter_029:sink0_startofpacket
	wire  [65:0] width_adapter_076_src_data;                                                              // width_adapter_076:out_data -> burst_adapter_029:sink0_data
	wire         width_adapter_076_src_ready;                                                             // burst_adapter_029:sink0_ready -> width_adapter_076:out_ready
	wire  [57:0] width_adapter_076_src_channel;                                                           // width_adapter_076:out_channel -> burst_adapter_029:sink0_channel
	wire         id_router_044_src_endofpacket;                                                           // id_router_044:src_endofpacket -> width_adapter_077:in_endofpacket
	wire         id_router_044_src_valid;                                                                 // id_router_044:src_valid -> width_adapter_077:in_valid
	wire         id_router_044_src_startofpacket;                                                         // id_router_044:src_startofpacket -> width_adapter_077:in_startofpacket
	wire  [65:0] id_router_044_src_data;                                                                  // id_router_044:src_data -> width_adapter_077:in_data
	wire  [57:0] id_router_044_src_channel;                                                               // id_router_044:src_channel -> width_adapter_077:in_channel
	wire         id_router_044_src_ready;                                                                 // width_adapter_077:in_ready -> id_router_044:src_ready
	wire         width_adapter_077_src_endofpacket;                                                       // width_adapter_077:out_endofpacket -> rsp_xbar_demux_044:sink_endofpacket
	wire         width_adapter_077_src_valid;                                                             // width_adapter_077:out_valid -> rsp_xbar_demux_044:sink_valid
	wire         width_adapter_077_src_startofpacket;                                                     // width_adapter_077:out_startofpacket -> rsp_xbar_demux_044:sink_startofpacket
	wire  [92:0] width_adapter_077_src_data;                                                              // width_adapter_077:out_data -> rsp_xbar_demux_044:sink_data
	wire         width_adapter_077_src_ready;                                                             // rsp_xbar_demux_044:sink_ready -> width_adapter_077:out_ready
	wire  [57:0] width_adapter_077_src_channel;                                                           // width_adapter_077:out_channel -> rsp_xbar_demux_044:sink_channel
	wire         cmd_xbar_demux_src45_ready;                                                              // width_adapter_078:in_ready -> cmd_xbar_demux:src45_ready
	wire         width_adapter_078_src_endofpacket;                                                       // width_adapter_078:out_endofpacket -> burst_adapter_035:sink0_endofpacket
	wire         width_adapter_078_src_valid;                                                             // width_adapter_078:out_valid -> burst_adapter_035:sink0_valid
	wire         width_adapter_078_src_startofpacket;                                                     // width_adapter_078:out_startofpacket -> burst_adapter_035:sink0_startofpacket
	wire  [65:0] width_adapter_078_src_data;                                                              // width_adapter_078:out_data -> burst_adapter_035:sink0_data
	wire         width_adapter_078_src_ready;                                                             // burst_adapter_035:sink0_ready -> width_adapter_078:out_ready
	wire  [57:0] width_adapter_078_src_channel;                                                           // width_adapter_078:out_channel -> burst_adapter_035:sink0_channel
	wire         id_router_045_src_endofpacket;                                                           // id_router_045:src_endofpacket -> width_adapter_079:in_endofpacket
	wire         id_router_045_src_valid;                                                                 // id_router_045:src_valid -> width_adapter_079:in_valid
	wire         id_router_045_src_startofpacket;                                                         // id_router_045:src_startofpacket -> width_adapter_079:in_startofpacket
	wire  [65:0] id_router_045_src_data;                                                                  // id_router_045:src_data -> width_adapter_079:in_data
	wire  [57:0] id_router_045_src_channel;                                                               // id_router_045:src_channel -> width_adapter_079:in_channel
	wire         id_router_045_src_ready;                                                                 // width_adapter_079:in_ready -> id_router_045:src_ready
	wire         width_adapter_079_src_endofpacket;                                                       // width_adapter_079:out_endofpacket -> rsp_xbar_demux_045:sink_endofpacket
	wire         width_adapter_079_src_valid;                                                             // width_adapter_079:out_valid -> rsp_xbar_demux_045:sink_valid
	wire         width_adapter_079_src_startofpacket;                                                     // width_adapter_079:out_startofpacket -> rsp_xbar_demux_045:sink_startofpacket
	wire  [92:0] width_adapter_079_src_data;                                                              // width_adapter_079:out_data -> rsp_xbar_demux_045:sink_data
	wire         width_adapter_079_src_ready;                                                             // rsp_xbar_demux_045:sink_ready -> width_adapter_079:out_ready
	wire  [57:0] width_adapter_079_src_channel;                                                           // width_adapter_079:out_channel -> rsp_xbar_demux_045:sink_channel
	wire         cmd_xbar_demux_src46_ready;                                                              // width_adapter_080:in_ready -> cmd_xbar_demux:src46_ready
	wire         width_adapter_080_src_endofpacket;                                                       // width_adapter_080:out_endofpacket -> burst_adapter_030:sink0_endofpacket
	wire         width_adapter_080_src_valid;                                                             // width_adapter_080:out_valid -> burst_adapter_030:sink0_valid
	wire         width_adapter_080_src_startofpacket;                                                     // width_adapter_080:out_startofpacket -> burst_adapter_030:sink0_startofpacket
	wire  [65:0] width_adapter_080_src_data;                                                              // width_adapter_080:out_data -> burst_adapter_030:sink0_data
	wire         width_adapter_080_src_ready;                                                             // burst_adapter_030:sink0_ready -> width_adapter_080:out_ready
	wire  [57:0] width_adapter_080_src_channel;                                                           // width_adapter_080:out_channel -> burst_adapter_030:sink0_channel
	wire         id_router_046_src_endofpacket;                                                           // id_router_046:src_endofpacket -> width_adapter_081:in_endofpacket
	wire         id_router_046_src_valid;                                                                 // id_router_046:src_valid -> width_adapter_081:in_valid
	wire         id_router_046_src_startofpacket;                                                         // id_router_046:src_startofpacket -> width_adapter_081:in_startofpacket
	wire  [65:0] id_router_046_src_data;                                                                  // id_router_046:src_data -> width_adapter_081:in_data
	wire  [57:0] id_router_046_src_channel;                                                               // id_router_046:src_channel -> width_adapter_081:in_channel
	wire         id_router_046_src_ready;                                                                 // width_adapter_081:in_ready -> id_router_046:src_ready
	wire         width_adapter_081_src_endofpacket;                                                       // width_adapter_081:out_endofpacket -> rsp_xbar_demux_046:sink_endofpacket
	wire         width_adapter_081_src_valid;                                                             // width_adapter_081:out_valid -> rsp_xbar_demux_046:sink_valid
	wire         width_adapter_081_src_startofpacket;                                                     // width_adapter_081:out_startofpacket -> rsp_xbar_demux_046:sink_startofpacket
	wire  [92:0] width_adapter_081_src_data;                                                              // width_adapter_081:out_data -> rsp_xbar_demux_046:sink_data
	wire         width_adapter_081_src_ready;                                                             // rsp_xbar_demux_046:sink_ready -> width_adapter_081:out_ready
	wire  [57:0] width_adapter_081_src_channel;                                                           // width_adapter_081:out_channel -> rsp_xbar_demux_046:sink_channel
	wire         cmd_xbar_demux_src47_ready;                                                              // width_adapter_082:in_ready -> cmd_xbar_demux:src47_ready
	wire         width_adapter_082_src_endofpacket;                                                       // width_adapter_082:out_endofpacket -> burst_adapter_022:sink0_endofpacket
	wire         width_adapter_082_src_valid;                                                             // width_adapter_082:out_valid -> burst_adapter_022:sink0_valid
	wire         width_adapter_082_src_startofpacket;                                                     // width_adapter_082:out_startofpacket -> burst_adapter_022:sink0_startofpacket
	wire  [65:0] width_adapter_082_src_data;                                                              // width_adapter_082:out_data -> burst_adapter_022:sink0_data
	wire         width_adapter_082_src_ready;                                                             // burst_adapter_022:sink0_ready -> width_adapter_082:out_ready
	wire  [57:0] width_adapter_082_src_channel;                                                           // width_adapter_082:out_channel -> burst_adapter_022:sink0_channel
	wire         id_router_047_src_endofpacket;                                                           // id_router_047:src_endofpacket -> width_adapter_083:in_endofpacket
	wire         id_router_047_src_valid;                                                                 // id_router_047:src_valid -> width_adapter_083:in_valid
	wire         id_router_047_src_startofpacket;                                                         // id_router_047:src_startofpacket -> width_adapter_083:in_startofpacket
	wire  [65:0] id_router_047_src_data;                                                                  // id_router_047:src_data -> width_adapter_083:in_data
	wire  [57:0] id_router_047_src_channel;                                                               // id_router_047:src_channel -> width_adapter_083:in_channel
	wire         id_router_047_src_ready;                                                                 // width_adapter_083:in_ready -> id_router_047:src_ready
	wire         width_adapter_083_src_endofpacket;                                                       // width_adapter_083:out_endofpacket -> rsp_xbar_demux_047:sink_endofpacket
	wire         width_adapter_083_src_valid;                                                             // width_adapter_083:out_valid -> rsp_xbar_demux_047:sink_valid
	wire         width_adapter_083_src_startofpacket;                                                     // width_adapter_083:out_startofpacket -> rsp_xbar_demux_047:sink_startofpacket
	wire  [92:0] width_adapter_083_src_data;                                                              // width_adapter_083:out_data -> rsp_xbar_demux_047:sink_data
	wire         width_adapter_083_src_ready;                                                             // rsp_xbar_demux_047:sink_ready -> width_adapter_083:out_ready
	wire  [57:0] width_adapter_083_src_channel;                                                           // width_adapter_083:out_channel -> rsp_xbar_demux_047:sink_channel
	wire         cmd_xbar_demux_src48_ready;                                                              // width_adapter_084:in_ready -> cmd_xbar_demux:src48_ready
	wire         width_adapter_084_src_endofpacket;                                                       // width_adapter_084:out_endofpacket -> burst_adapter_020:sink0_endofpacket
	wire         width_adapter_084_src_valid;                                                             // width_adapter_084:out_valid -> burst_adapter_020:sink0_valid
	wire         width_adapter_084_src_startofpacket;                                                     // width_adapter_084:out_startofpacket -> burst_adapter_020:sink0_startofpacket
	wire  [65:0] width_adapter_084_src_data;                                                              // width_adapter_084:out_data -> burst_adapter_020:sink0_data
	wire         width_adapter_084_src_ready;                                                             // burst_adapter_020:sink0_ready -> width_adapter_084:out_ready
	wire  [57:0] width_adapter_084_src_channel;                                                           // width_adapter_084:out_channel -> burst_adapter_020:sink0_channel
	wire         id_router_048_src_endofpacket;                                                           // id_router_048:src_endofpacket -> width_adapter_085:in_endofpacket
	wire         id_router_048_src_valid;                                                                 // id_router_048:src_valid -> width_adapter_085:in_valid
	wire         id_router_048_src_startofpacket;                                                         // id_router_048:src_startofpacket -> width_adapter_085:in_startofpacket
	wire  [65:0] id_router_048_src_data;                                                                  // id_router_048:src_data -> width_adapter_085:in_data
	wire  [57:0] id_router_048_src_channel;                                                               // id_router_048:src_channel -> width_adapter_085:in_channel
	wire         id_router_048_src_ready;                                                                 // width_adapter_085:in_ready -> id_router_048:src_ready
	wire         width_adapter_085_src_endofpacket;                                                       // width_adapter_085:out_endofpacket -> rsp_xbar_demux_048:sink_endofpacket
	wire         width_adapter_085_src_valid;                                                             // width_adapter_085:out_valid -> rsp_xbar_demux_048:sink_valid
	wire         width_adapter_085_src_startofpacket;                                                     // width_adapter_085:out_startofpacket -> rsp_xbar_demux_048:sink_startofpacket
	wire  [92:0] width_adapter_085_src_data;                                                              // width_adapter_085:out_data -> rsp_xbar_demux_048:sink_data
	wire         width_adapter_085_src_ready;                                                             // rsp_xbar_demux_048:sink_ready -> width_adapter_085:out_ready
	wire  [57:0] width_adapter_085_src_channel;                                                           // width_adapter_085:out_channel -> rsp_xbar_demux_048:sink_channel
	wire         cmd_xbar_demux_src49_ready;                                                              // width_adapter_086:in_ready -> cmd_xbar_demux:src49_ready
	wire         width_adapter_086_src_endofpacket;                                                       // width_adapter_086:out_endofpacket -> burst_adapter_045:sink0_endofpacket
	wire         width_adapter_086_src_valid;                                                             // width_adapter_086:out_valid -> burst_adapter_045:sink0_valid
	wire         width_adapter_086_src_startofpacket;                                                     // width_adapter_086:out_startofpacket -> burst_adapter_045:sink0_startofpacket
	wire  [65:0] width_adapter_086_src_data;                                                              // width_adapter_086:out_data -> burst_adapter_045:sink0_data
	wire         width_adapter_086_src_ready;                                                             // burst_adapter_045:sink0_ready -> width_adapter_086:out_ready
	wire  [57:0] width_adapter_086_src_channel;                                                           // width_adapter_086:out_channel -> burst_adapter_045:sink0_channel
	wire         id_router_049_src_endofpacket;                                                           // id_router_049:src_endofpacket -> width_adapter_087:in_endofpacket
	wire         id_router_049_src_valid;                                                                 // id_router_049:src_valid -> width_adapter_087:in_valid
	wire         id_router_049_src_startofpacket;                                                         // id_router_049:src_startofpacket -> width_adapter_087:in_startofpacket
	wire  [65:0] id_router_049_src_data;                                                                  // id_router_049:src_data -> width_adapter_087:in_data
	wire  [57:0] id_router_049_src_channel;                                                               // id_router_049:src_channel -> width_adapter_087:in_channel
	wire         id_router_049_src_ready;                                                                 // width_adapter_087:in_ready -> id_router_049:src_ready
	wire         width_adapter_087_src_endofpacket;                                                       // width_adapter_087:out_endofpacket -> rsp_xbar_demux_049:sink_endofpacket
	wire         width_adapter_087_src_valid;                                                             // width_adapter_087:out_valid -> rsp_xbar_demux_049:sink_valid
	wire         width_adapter_087_src_startofpacket;                                                     // width_adapter_087:out_startofpacket -> rsp_xbar_demux_049:sink_startofpacket
	wire  [92:0] width_adapter_087_src_data;                                                              // width_adapter_087:out_data -> rsp_xbar_demux_049:sink_data
	wire         width_adapter_087_src_ready;                                                             // rsp_xbar_demux_049:sink_ready -> width_adapter_087:out_ready
	wire  [57:0] width_adapter_087_src_channel;                                                           // width_adapter_087:out_channel -> rsp_xbar_demux_049:sink_channel
	wire         cmd_xbar_demux_src50_ready;                                                              // width_adapter_088:in_ready -> cmd_xbar_demux:src50_ready
	wire         width_adapter_088_src_endofpacket;                                                       // width_adapter_088:out_endofpacket -> burst_adapter_038:sink0_endofpacket
	wire         width_adapter_088_src_valid;                                                             // width_adapter_088:out_valid -> burst_adapter_038:sink0_valid
	wire         width_adapter_088_src_startofpacket;                                                     // width_adapter_088:out_startofpacket -> burst_adapter_038:sink0_startofpacket
	wire  [65:0] width_adapter_088_src_data;                                                              // width_adapter_088:out_data -> burst_adapter_038:sink0_data
	wire         width_adapter_088_src_ready;                                                             // burst_adapter_038:sink0_ready -> width_adapter_088:out_ready
	wire  [57:0] width_adapter_088_src_channel;                                                           // width_adapter_088:out_channel -> burst_adapter_038:sink0_channel
	wire         id_router_050_src_endofpacket;                                                           // id_router_050:src_endofpacket -> width_adapter_089:in_endofpacket
	wire         id_router_050_src_valid;                                                                 // id_router_050:src_valid -> width_adapter_089:in_valid
	wire         id_router_050_src_startofpacket;                                                         // id_router_050:src_startofpacket -> width_adapter_089:in_startofpacket
	wire  [65:0] id_router_050_src_data;                                                                  // id_router_050:src_data -> width_adapter_089:in_data
	wire  [57:0] id_router_050_src_channel;                                                               // id_router_050:src_channel -> width_adapter_089:in_channel
	wire         id_router_050_src_ready;                                                                 // width_adapter_089:in_ready -> id_router_050:src_ready
	wire         width_adapter_089_src_endofpacket;                                                       // width_adapter_089:out_endofpacket -> rsp_xbar_demux_050:sink_endofpacket
	wire         width_adapter_089_src_valid;                                                             // width_adapter_089:out_valid -> rsp_xbar_demux_050:sink_valid
	wire         width_adapter_089_src_startofpacket;                                                     // width_adapter_089:out_startofpacket -> rsp_xbar_demux_050:sink_startofpacket
	wire  [92:0] width_adapter_089_src_data;                                                              // width_adapter_089:out_data -> rsp_xbar_demux_050:sink_data
	wire         width_adapter_089_src_ready;                                                             // rsp_xbar_demux_050:sink_ready -> width_adapter_089:out_ready
	wire  [57:0] width_adapter_089_src_channel;                                                           // width_adapter_089:out_channel -> rsp_xbar_demux_050:sink_channel
	wire         cmd_xbar_demux_src51_ready;                                                              // width_adapter_090:in_ready -> cmd_xbar_demux:src51_ready
	wire         width_adapter_090_src_endofpacket;                                                       // width_adapter_090:out_endofpacket -> burst_adapter_006:sink0_endofpacket
	wire         width_adapter_090_src_valid;                                                             // width_adapter_090:out_valid -> burst_adapter_006:sink0_valid
	wire         width_adapter_090_src_startofpacket;                                                     // width_adapter_090:out_startofpacket -> burst_adapter_006:sink0_startofpacket
	wire  [65:0] width_adapter_090_src_data;                                                              // width_adapter_090:out_data -> burst_adapter_006:sink0_data
	wire         width_adapter_090_src_ready;                                                             // burst_adapter_006:sink0_ready -> width_adapter_090:out_ready
	wire  [57:0] width_adapter_090_src_channel;                                                           // width_adapter_090:out_channel -> burst_adapter_006:sink0_channel
	wire         id_router_051_src_endofpacket;                                                           // id_router_051:src_endofpacket -> width_adapter_091:in_endofpacket
	wire         id_router_051_src_valid;                                                                 // id_router_051:src_valid -> width_adapter_091:in_valid
	wire         id_router_051_src_startofpacket;                                                         // id_router_051:src_startofpacket -> width_adapter_091:in_startofpacket
	wire  [65:0] id_router_051_src_data;                                                                  // id_router_051:src_data -> width_adapter_091:in_data
	wire  [57:0] id_router_051_src_channel;                                                               // id_router_051:src_channel -> width_adapter_091:in_channel
	wire         id_router_051_src_ready;                                                                 // width_adapter_091:in_ready -> id_router_051:src_ready
	wire         width_adapter_091_src_endofpacket;                                                       // width_adapter_091:out_endofpacket -> rsp_xbar_demux_051:sink_endofpacket
	wire         width_adapter_091_src_valid;                                                             // width_adapter_091:out_valid -> rsp_xbar_demux_051:sink_valid
	wire         width_adapter_091_src_startofpacket;                                                     // width_adapter_091:out_startofpacket -> rsp_xbar_demux_051:sink_startofpacket
	wire  [92:0] width_adapter_091_src_data;                                                              // width_adapter_091:out_data -> rsp_xbar_demux_051:sink_data
	wire         width_adapter_091_src_ready;                                                             // rsp_xbar_demux_051:sink_ready -> width_adapter_091:out_ready
	wire  [57:0] width_adapter_091_src_channel;                                                           // width_adapter_091:out_channel -> rsp_xbar_demux_051:sink_channel
	wire         cmd_xbar_demux_src52_ready;                                                              // width_adapter_092:in_ready -> cmd_xbar_demux:src52_ready
	wire         width_adapter_092_src_endofpacket;                                                       // width_adapter_092:out_endofpacket -> burst_adapter_018:sink0_endofpacket
	wire         width_adapter_092_src_valid;                                                             // width_adapter_092:out_valid -> burst_adapter_018:sink0_valid
	wire         width_adapter_092_src_startofpacket;                                                     // width_adapter_092:out_startofpacket -> burst_adapter_018:sink0_startofpacket
	wire  [65:0] width_adapter_092_src_data;                                                              // width_adapter_092:out_data -> burst_adapter_018:sink0_data
	wire         width_adapter_092_src_ready;                                                             // burst_adapter_018:sink0_ready -> width_adapter_092:out_ready
	wire  [57:0] width_adapter_092_src_channel;                                                           // width_adapter_092:out_channel -> burst_adapter_018:sink0_channel
	wire         id_router_052_src_endofpacket;                                                           // id_router_052:src_endofpacket -> width_adapter_093:in_endofpacket
	wire         id_router_052_src_valid;                                                                 // id_router_052:src_valid -> width_adapter_093:in_valid
	wire         id_router_052_src_startofpacket;                                                         // id_router_052:src_startofpacket -> width_adapter_093:in_startofpacket
	wire  [65:0] id_router_052_src_data;                                                                  // id_router_052:src_data -> width_adapter_093:in_data
	wire  [57:0] id_router_052_src_channel;                                                               // id_router_052:src_channel -> width_adapter_093:in_channel
	wire         id_router_052_src_ready;                                                                 // width_adapter_093:in_ready -> id_router_052:src_ready
	wire         width_adapter_093_src_endofpacket;                                                       // width_adapter_093:out_endofpacket -> rsp_xbar_demux_052:sink_endofpacket
	wire         width_adapter_093_src_valid;                                                             // width_adapter_093:out_valid -> rsp_xbar_demux_052:sink_valid
	wire         width_adapter_093_src_startofpacket;                                                     // width_adapter_093:out_startofpacket -> rsp_xbar_demux_052:sink_startofpacket
	wire  [92:0] width_adapter_093_src_data;                                                              // width_adapter_093:out_data -> rsp_xbar_demux_052:sink_data
	wire         width_adapter_093_src_ready;                                                             // rsp_xbar_demux_052:sink_ready -> width_adapter_093:out_ready
	wire  [57:0] width_adapter_093_src_channel;                                                           // width_adapter_093:out_channel -> rsp_xbar_demux_052:sink_channel
	wire         cmd_xbar_demux_src53_ready;                                                              // width_adapter_094:in_ready -> cmd_xbar_demux:src53_ready
	wire         width_adapter_094_src_endofpacket;                                                       // width_adapter_094:out_endofpacket -> burst_adapter_024:sink0_endofpacket
	wire         width_adapter_094_src_valid;                                                             // width_adapter_094:out_valid -> burst_adapter_024:sink0_valid
	wire         width_adapter_094_src_startofpacket;                                                     // width_adapter_094:out_startofpacket -> burst_adapter_024:sink0_startofpacket
	wire  [65:0] width_adapter_094_src_data;                                                              // width_adapter_094:out_data -> burst_adapter_024:sink0_data
	wire         width_adapter_094_src_ready;                                                             // burst_adapter_024:sink0_ready -> width_adapter_094:out_ready
	wire  [57:0] width_adapter_094_src_channel;                                                           // width_adapter_094:out_channel -> burst_adapter_024:sink0_channel
	wire         id_router_053_src_endofpacket;                                                           // id_router_053:src_endofpacket -> width_adapter_095:in_endofpacket
	wire         id_router_053_src_valid;                                                                 // id_router_053:src_valid -> width_adapter_095:in_valid
	wire         id_router_053_src_startofpacket;                                                         // id_router_053:src_startofpacket -> width_adapter_095:in_startofpacket
	wire  [65:0] id_router_053_src_data;                                                                  // id_router_053:src_data -> width_adapter_095:in_data
	wire  [57:0] id_router_053_src_channel;                                                               // id_router_053:src_channel -> width_adapter_095:in_channel
	wire         id_router_053_src_ready;                                                                 // width_adapter_095:in_ready -> id_router_053:src_ready
	wire         width_adapter_095_src_endofpacket;                                                       // width_adapter_095:out_endofpacket -> rsp_xbar_demux_053:sink_endofpacket
	wire         width_adapter_095_src_valid;                                                             // width_adapter_095:out_valid -> rsp_xbar_demux_053:sink_valid
	wire         width_adapter_095_src_startofpacket;                                                     // width_adapter_095:out_startofpacket -> rsp_xbar_demux_053:sink_startofpacket
	wire  [92:0] width_adapter_095_src_data;                                                              // width_adapter_095:out_data -> rsp_xbar_demux_053:sink_data
	wire         width_adapter_095_src_ready;                                                             // rsp_xbar_demux_053:sink_ready -> width_adapter_095:out_ready
	wire  [57:0] width_adapter_095_src_channel;                                                           // width_adapter_095:out_channel -> rsp_xbar_demux_053:sink_channel
	wire         cmd_xbar_demux_src54_ready;                                                              // width_adapter_096:in_ready -> cmd_xbar_demux:src54_ready
	wire         width_adapter_096_src_endofpacket;                                                       // width_adapter_096:out_endofpacket -> burst_adapter_039:sink0_endofpacket
	wire         width_adapter_096_src_valid;                                                             // width_adapter_096:out_valid -> burst_adapter_039:sink0_valid
	wire         width_adapter_096_src_startofpacket;                                                     // width_adapter_096:out_startofpacket -> burst_adapter_039:sink0_startofpacket
	wire  [65:0] width_adapter_096_src_data;                                                              // width_adapter_096:out_data -> burst_adapter_039:sink0_data
	wire         width_adapter_096_src_ready;                                                             // burst_adapter_039:sink0_ready -> width_adapter_096:out_ready
	wire  [57:0] width_adapter_096_src_channel;                                                           // width_adapter_096:out_channel -> burst_adapter_039:sink0_channel
	wire         id_router_054_src_endofpacket;                                                           // id_router_054:src_endofpacket -> width_adapter_097:in_endofpacket
	wire         id_router_054_src_valid;                                                                 // id_router_054:src_valid -> width_adapter_097:in_valid
	wire         id_router_054_src_startofpacket;                                                         // id_router_054:src_startofpacket -> width_adapter_097:in_startofpacket
	wire  [65:0] id_router_054_src_data;                                                                  // id_router_054:src_data -> width_adapter_097:in_data
	wire  [57:0] id_router_054_src_channel;                                                               // id_router_054:src_channel -> width_adapter_097:in_channel
	wire         id_router_054_src_ready;                                                                 // width_adapter_097:in_ready -> id_router_054:src_ready
	wire         width_adapter_097_src_endofpacket;                                                       // width_adapter_097:out_endofpacket -> rsp_xbar_demux_054:sink_endofpacket
	wire         width_adapter_097_src_valid;                                                             // width_adapter_097:out_valid -> rsp_xbar_demux_054:sink_valid
	wire         width_adapter_097_src_startofpacket;                                                     // width_adapter_097:out_startofpacket -> rsp_xbar_demux_054:sink_startofpacket
	wire  [92:0] width_adapter_097_src_data;                                                              // width_adapter_097:out_data -> rsp_xbar_demux_054:sink_data
	wire         width_adapter_097_src_ready;                                                             // rsp_xbar_demux_054:sink_ready -> width_adapter_097:out_ready
	wire  [57:0] width_adapter_097_src_channel;                                                           // width_adapter_097:out_channel -> rsp_xbar_demux_054:sink_channel
	wire         cmd_xbar_demux_src55_ready;                                                              // width_adapter_098:in_ready -> cmd_xbar_demux:src55_ready
	wire         width_adapter_098_src_endofpacket;                                                       // width_adapter_098:out_endofpacket -> burst_adapter_034:sink0_endofpacket
	wire         width_adapter_098_src_valid;                                                             // width_adapter_098:out_valid -> burst_adapter_034:sink0_valid
	wire         width_adapter_098_src_startofpacket;                                                     // width_adapter_098:out_startofpacket -> burst_adapter_034:sink0_startofpacket
	wire  [65:0] width_adapter_098_src_data;                                                              // width_adapter_098:out_data -> burst_adapter_034:sink0_data
	wire         width_adapter_098_src_ready;                                                             // burst_adapter_034:sink0_ready -> width_adapter_098:out_ready
	wire  [57:0] width_adapter_098_src_channel;                                                           // width_adapter_098:out_channel -> burst_adapter_034:sink0_channel
	wire         id_router_055_src_endofpacket;                                                           // id_router_055:src_endofpacket -> width_adapter_099:in_endofpacket
	wire         id_router_055_src_valid;                                                                 // id_router_055:src_valid -> width_adapter_099:in_valid
	wire         id_router_055_src_startofpacket;                                                         // id_router_055:src_startofpacket -> width_adapter_099:in_startofpacket
	wire  [65:0] id_router_055_src_data;                                                                  // id_router_055:src_data -> width_adapter_099:in_data
	wire  [57:0] id_router_055_src_channel;                                                               // id_router_055:src_channel -> width_adapter_099:in_channel
	wire         id_router_055_src_ready;                                                                 // width_adapter_099:in_ready -> id_router_055:src_ready
	wire         width_adapter_099_src_endofpacket;                                                       // width_adapter_099:out_endofpacket -> rsp_xbar_demux_055:sink_endofpacket
	wire         width_adapter_099_src_valid;                                                             // width_adapter_099:out_valid -> rsp_xbar_demux_055:sink_valid
	wire         width_adapter_099_src_startofpacket;                                                     // width_adapter_099:out_startofpacket -> rsp_xbar_demux_055:sink_startofpacket
	wire  [92:0] width_adapter_099_src_data;                                                              // width_adapter_099:out_data -> rsp_xbar_demux_055:sink_data
	wire         width_adapter_099_src_ready;                                                             // rsp_xbar_demux_055:sink_ready -> width_adapter_099:out_ready
	wire  [57:0] width_adapter_099_src_channel;                                                           // width_adapter_099:out_channel -> rsp_xbar_demux_055:sink_channel
	wire         cmd_xbar_demux_src56_ready;                                                              // width_adapter_100:in_ready -> cmd_xbar_demux:src56_ready
	wire         width_adapter_100_src_endofpacket;                                                       // width_adapter_100:out_endofpacket -> burst_adapter_016:sink0_endofpacket
	wire         width_adapter_100_src_valid;                                                             // width_adapter_100:out_valid -> burst_adapter_016:sink0_valid
	wire         width_adapter_100_src_startofpacket;                                                     // width_adapter_100:out_startofpacket -> burst_adapter_016:sink0_startofpacket
	wire  [65:0] width_adapter_100_src_data;                                                              // width_adapter_100:out_data -> burst_adapter_016:sink0_data
	wire         width_adapter_100_src_ready;                                                             // burst_adapter_016:sink0_ready -> width_adapter_100:out_ready
	wire  [57:0] width_adapter_100_src_channel;                                                           // width_adapter_100:out_channel -> burst_adapter_016:sink0_channel
	wire         id_router_056_src_endofpacket;                                                           // id_router_056:src_endofpacket -> width_adapter_101:in_endofpacket
	wire         id_router_056_src_valid;                                                                 // id_router_056:src_valid -> width_adapter_101:in_valid
	wire         id_router_056_src_startofpacket;                                                         // id_router_056:src_startofpacket -> width_adapter_101:in_startofpacket
	wire  [65:0] id_router_056_src_data;                                                                  // id_router_056:src_data -> width_adapter_101:in_data
	wire  [57:0] id_router_056_src_channel;                                                               // id_router_056:src_channel -> width_adapter_101:in_channel
	wire         id_router_056_src_ready;                                                                 // width_adapter_101:in_ready -> id_router_056:src_ready
	wire         width_adapter_101_src_endofpacket;                                                       // width_adapter_101:out_endofpacket -> rsp_xbar_demux_056:sink_endofpacket
	wire         width_adapter_101_src_valid;                                                             // width_adapter_101:out_valid -> rsp_xbar_demux_056:sink_valid
	wire         width_adapter_101_src_startofpacket;                                                     // width_adapter_101:out_startofpacket -> rsp_xbar_demux_056:sink_startofpacket
	wire  [92:0] width_adapter_101_src_data;                                                              // width_adapter_101:out_data -> rsp_xbar_demux_056:sink_data
	wire         width_adapter_101_src_ready;                                                             // rsp_xbar_demux_056:sink_ready -> width_adapter_101:out_ready
	wire  [57:0] width_adapter_101_src_channel;                                                           // width_adapter_101:out_channel -> rsp_xbar_demux_056:sink_channel
	wire         cmd_xbar_demux_src57_ready;                                                              // width_adapter_102:in_ready -> cmd_xbar_demux:src57_ready
	wire         width_adapter_102_src_endofpacket;                                                       // width_adapter_102:out_endofpacket -> burst_adapter_036:sink0_endofpacket
	wire         width_adapter_102_src_valid;                                                             // width_adapter_102:out_valid -> burst_adapter_036:sink0_valid
	wire         width_adapter_102_src_startofpacket;                                                     // width_adapter_102:out_startofpacket -> burst_adapter_036:sink0_startofpacket
	wire  [65:0] width_adapter_102_src_data;                                                              // width_adapter_102:out_data -> burst_adapter_036:sink0_data
	wire         width_adapter_102_src_ready;                                                             // burst_adapter_036:sink0_ready -> width_adapter_102:out_ready
	wire  [57:0] width_adapter_102_src_channel;                                                           // width_adapter_102:out_channel -> burst_adapter_036:sink0_channel
	wire         id_router_057_src_endofpacket;                                                           // id_router_057:src_endofpacket -> width_adapter_103:in_endofpacket
	wire         id_router_057_src_valid;                                                                 // id_router_057:src_valid -> width_adapter_103:in_valid
	wire         id_router_057_src_startofpacket;                                                         // id_router_057:src_startofpacket -> width_adapter_103:in_startofpacket
	wire  [65:0] id_router_057_src_data;                                                                  // id_router_057:src_data -> width_adapter_103:in_data
	wire  [57:0] id_router_057_src_channel;                                                               // id_router_057:src_channel -> width_adapter_103:in_channel
	wire         id_router_057_src_ready;                                                                 // width_adapter_103:in_ready -> id_router_057:src_ready
	wire         width_adapter_103_src_endofpacket;                                                       // width_adapter_103:out_endofpacket -> rsp_xbar_demux_057:sink_endofpacket
	wire         width_adapter_103_src_valid;                                                             // width_adapter_103:out_valid -> rsp_xbar_demux_057:sink_valid
	wire         width_adapter_103_src_startofpacket;                                                     // width_adapter_103:out_startofpacket -> rsp_xbar_demux_057:sink_startofpacket
	wire  [92:0] width_adapter_103_src_data;                                                              // width_adapter_103:out_data -> rsp_xbar_demux_057:sink_data
	wire         width_adapter_103_src_ready;                                                             // rsp_xbar_demux_057:sink_ready -> width_adapter_103:out_ready
	wire  [57:0] width_adapter_103_src_channel;                                                           // width_adapter_103:out_channel -> rsp_xbar_demux_057:sink_channel
	wire  [57:0] limiter_cmd_valid_data;                                                                  // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                // Shield_Admin:ins_OC_irq -> irq_mapper:receiver0_irq
	wire   [9:0] sam9_events_irq;                                                                         // irq_synchronizer:sender_irq -> SAM9:inr_EVENTS_irq
	wire   [9:0] irq_synchronizer_receiver_irq;                                                           // irq_mapper:sender_irq -> irq_synchronizer:receiver_irq

	qsys_tabby_host sam9 (
		.rso_MRST_reset       (sam9_mrst_reset),       //   MRST.reset
		.cso_MCLK_clk         (sam9_mclk_clk),         //   MCLK.clk
		.cso_H1CLK_clk        (),                      //  H1CLK.clk
		.cso_H2CLK_clk        (),                      //  H2CLK.clk
		.avm_M1_writedata     (sam9_m1_writedata),     //     M1.writedata
		.avm_M1_readdata      (sam9_m1_readdata),      //       .readdata
		.avm_M1_address       (sam9_m1_address),       //       .address
		.avm_M1_byteenable    (sam9_m1_byteenable),    //       .byteenable
		.avm_M1_write         (sam9_m1_write),         //       .write
		.avm_M1_read          (sam9_m1_read),          //       .read
		.avm_M1_begintransfer (sam9_m1_begintransfer), //       .begintransfer
		.avm_M1_readdatavalid (sam9_m1_readdatavalid), //       .readdatavalid
		.avm_M1_waitrequest   (sam9_m1_waitrequest),   //       .waitrequest
		.inr_EVENTS_irq       (sam9_events_irq),       // EVENTS.irq
		.coe_M1_RSTN          (m1_RSTN),               // EXPORT.export
		.coe_M1_CLK           (m1_CLK),                //       .export
		.coe_M1_ADDR          (m1_ADDR),               //       .export
		.coe_M1_DATA          (m1_DATA),               //       .export
		.coe_M1_CSN           (m1_CSN),                //       .export
		.coe_M1_BEN           (m1_BEN),                //       .export
		.coe_M1_RDN           (m1_RDN),                //       .export
		.coe_M1_WRN           (m1_WRN),                //       .export
		.coe_M1_WAITN         (m1_WAITN),              //       .export
		.coe_M1_EINT          (m1_EINT)                //       .export
	);

	qsys_basic_SysID sysid (
		.rsi_MRST_reset        (sam9_mrst_reset),                                        //  MRST.reset
		.csi_MCLK_clk          (sam9_mclk_clk),                                          //  MCLK.clk
		.avs_SysID_readdata    (sysid_sysid_translator_avalon_anti_slave_0_readdata),    // SysID.readdata
		.avs_SysID_read        (sysid_sysid_translator_avalon_anti_slave_0_read),        //      .read
		.avs_SysID_waitrequest (sysid_sysid_translator_avalon_anti_slave_0_waitrequest)  //      .waitrequest
	);

	qsys_basic_FuncLED funcled_0 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                           //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                             //   MCLK.clk
		.avs_LEDD_writedata   (funcled_0_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (funcled_0_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (funcled_0_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (funcled_0_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (funcled_0_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (funcled_0_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (qsys_test_ledstate_0_leds_data),                            //   LEDS.data
		.asi_LEDS_valid       (qsys_test_ledstate_0_leds_valid),                           //       .valid
		.asi_LEDS_ready       (qsys_test_ledstate_0_leds_ready),                           //       .ready
		.coe_LED_R            (led_f0_R),                                                  // EXPORT.export
		.coe_LED_G            (led_f0_G),                                                  //       .export
		.coe_LED_B            (led_f0_B)                                                   //       .export
	);

	qsys_basic_FuncLED funcled_1 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                           //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                             //   MCLK.clk
		.avs_LEDD_writedata   (funcled_1_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (funcled_1_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (funcled_1_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (funcled_1_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (funcled_1_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (funcled_1_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (qsys_test_ledstate_1_leds_data),                            //   LEDS.data
		.asi_LEDS_valid       (qsys_test_ledstate_1_leds_valid),                           //       .valid
		.asi_LEDS_ready       (qsys_test_ledstate_1_leds_ready),                           //       .ready
		.coe_LED_R            (led_f1_R),                                                  // EXPORT.export
		.coe_LED_G            (led_f1_G),                                                  //       .export
		.coe_LED_B            (led_f1_B)                                                   //       .export
	);

	qsys_basic_FuncLED funcled_2 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                           //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                             //   MCLK.clk
		.avs_LEDD_writedata   (funcled_2_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (funcled_2_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (funcled_2_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (funcled_2_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (funcled_2_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (funcled_2_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (qsys_test_ledstate_2_leds_data),                            //   LEDS.data
		.asi_LEDS_valid       (qsys_test_ledstate_2_leds_valid),                           //       .valid
		.asi_LEDS_ready       (qsys_test_ledstate_2_leds_ready),                           //       .ready
		.coe_LED_R            (led_f2_R),                                                  // EXPORT.export
		.coe_LED_G            (led_f2_G),                                                  //       .export
		.coe_LED_B            (led_f2_B)                                                   //       .export
	);

	qsys_basic_FuncLED funcled_3 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                           //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                             //   MCLK.clk
		.avs_LEDD_writedata   (funcled_3_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (funcled_3_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (funcled_3_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (funcled_3_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (funcled_3_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (funcled_3_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (qsys_test_ledstate_3_leds_data),                            //   LEDS.data
		.asi_LEDS_valid       (qsys_test_ledstate_3_leds_valid),                           //       .valid
		.asi_LEDS_ready       (qsys_test_ledstate_3_leds_ready),                           //       .ready
		.coe_LED_R            (led_f3_R),                                                  // EXPORT.export
		.coe_LED_G            (led_f3_G),                                                  //       .export
		.coe_LED_B            (led_f3_B)                                                   //       .export
	);

	qsys_shield_moduleBasicCtrl shield_admin (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_Ctrl_writedata   (shield_admin_ctrl_translator_avalon_anti_slave_0_writedata),   //   Ctrl.writedata
		.avs_Ctrl_readdata    (shield_admin_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_Ctrl_byteenable  (shield_admin_ctrl_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_Ctrl_write       (shield_admin_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_Ctrl_read        (shield_admin_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_Ctrl_waitrequest (shield_admin_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.ins_OC_irq           (irq_mapper_receiver0_irq),                                     //     OC.irq
		.coe_A_OCN            (shield_A_OCN),                                                 // EXPORT.export
		.coe_A_PWREN          (shield_A_PWREN),                                               //       .export
		.coe_A_HOE            (shield_A_HOE),                                                 //       .export
		.coe_A_LOE            (shield_A_LOE),                                                 //       .export
		.coe_B_OCN            (shield_B_OCN),                                                 //       .export
		.coe_B_PWREN          (shield_B_PWREN),                                               //       .export
		.coe_B_HOE            (shield_B_HOE),                                                 //       .export
		.coe_B_LOE            (shield_B_LOE)                                                  //       .export
	);

	qsys_test_LEDState qsys_test_ledstate_0 (
		.rsi_MRST_reset (sam9_mrst_reset),                 // MRST.reset
		.csi_MCLK_clk   (sam9_mclk_clk),                   // MCLK.clk
		.aso_LEDS_data  (qsys_test_ledstate_0_leds_data),  // LEDS.data
		.aso_LEDS_valid (qsys_test_ledstate_0_leds_valid), //     .valid
		.aso_LEDS_ready (qsys_test_ledstate_0_leds_ready)  //     .ready
	);

	qsys_test_LEDState qsys_test_ledstate_1 (
		.rsi_MRST_reset (sam9_mrst_reset),                 // MRST.reset
		.csi_MCLK_clk   (sam9_mclk_clk),                   // MCLK.clk
		.aso_LEDS_data  (qsys_test_ledstate_1_leds_data),  // LEDS.data
		.aso_LEDS_valid (qsys_test_ledstate_1_leds_valid), //     .valid
		.aso_LEDS_ready (qsys_test_ledstate_1_leds_ready)  //     .ready
	);

	qsys_test_LEDState qsys_test_ledstate_2 (
		.rsi_MRST_reset (sam9_mrst_reset),                 // MRST.reset
		.csi_MCLK_clk   (sam9_mclk_clk),                   // MCLK.clk
		.aso_LEDS_data  (qsys_test_ledstate_2_leds_data),  // LEDS.data
		.aso_LEDS_valid (qsys_test_ledstate_2_leds_valid), //     .valid
		.aso_LEDS_ready (qsys_test_ledstate_2_leds_ready)  //     .ready
	);

	qsys_test_LEDState qsys_test_ledstate_3 (
		.rsi_MRST_reset (sam9_mrst_reset),                 // MRST.reset
		.csi_MCLK_clk   (sam9_mclk_clk),                   // MCLK.clk
		.aso_LEDS_data  (qsys_test_ledstate_3_leds_data),  // LEDS.data
		.aso_LEDS_valid (qsys_test_ledstate_3_leds_valid), //     .valid
		.aso_LEDS_ready (qsys_test_ledstate_3_leds_ready)  //     .ready
	);

	qsys_shield_gpioFuncSel shiled_io_a0 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a0_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a0_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a0_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a0_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a0_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a0_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a0_f1_oe),                                                     //       .export
		.coe_f2_oe            (a0_f2_oe),                                                     //       .export
		.coe_f3_oe            (a0_f3_oe),                                                     //       .export
		.coe_f4_oe            (a0_f4_oe),                                                     //       .export
		.coe_f5_oe            (a0_f5_oe),                                                     //       .export
		.coe_f6_oe            (a0_f6_oe),                                                     //       .export
		.coe_f7_oe            (a0_f7_oe),                                                     //       .export
		.coe_f0_out           (a0_f0_out),                                                    //       .export
		.coe_f1_out           (a0_f1_out),                                                    //       .export
		.coe_f2_out           (a0_f2_out),                                                    //       .export
		.coe_f3_out           (a0_f3_out),                                                    //       .export
		.coe_f4_out           (a0_f4_out),                                                    //       .export
		.coe_f5_out           (a0_f5_out),                                                    //       .export
		.coe_f6_out           (a0_f6_out),                                                    //       .export
		.coe_f7_out           (a0_f7_out),                                                    //       .export
		.coe_f_in             (a0_f_in),                                                      //       .export
		.coe_GPIO             (a0_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a1 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a1_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a1_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a1_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a1_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a1_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a1_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a1_f1_oe),                                                     //       .export
		.coe_f2_oe            (a1_f2_oe),                                                     //       .export
		.coe_f3_oe            (a1_f3_oe),                                                     //       .export
		.coe_f4_oe            (a1_f4_oe),                                                     //       .export
		.coe_f5_oe            (a1_f5_oe),                                                     //       .export
		.coe_f6_oe            (a1_f6_oe),                                                     //       .export
		.coe_f7_oe            (a1_f7_oe),                                                     //       .export
		.coe_f0_out           (a1_f0_out),                                                    //       .export
		.coe_f1_out           (a1_f1_out),                                                    //       .export
		.coe_f2_out           (a1_f2_out),                                                    //       .export
		.coe_f3_out           (a1_f3_out),                                                    //       .export
		.coe_f4_out           (a1_f4_out),                                                    //       .export
		.coe_f5_out           (a1_f5_out),                                                    //       .export
		.coe_f6_out           (a1_f6_out),                                                    //       .export
		.coe_f7_out           (a1_f7_out),                                                    //       .export
		.coe_f_in             (a1_f_in),                                                      //       .export
		.coe_GPIO             (a1_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a2 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a2_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a2_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a2_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a2_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a2_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a2_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a2_f1_oe),                                                     //       .export
		.coe_f2_oe            (a2_f2_oe),                                                     //       .export
		.coe_f3_oe            (a2_f3_oe),                                                     //       .export
		.coe_f4_oe            (a2_f4_oe),                                                     //       .export
		.coe_f5_oe            (a2_f5_oe),                                                     //       .export
		.coe_f6_oe            (a2_f6_oe),                                                     //       .export
		.coe_f7_oe            (a2_f7_oe),                                                     //       .export
		.coe_f0_out           (a2_f0_out),                                                    //       .export
		.coe_f1_out           (a2_f1_out),                                                    //       .export
		.coe_f2_out           (a2_f2_out),                                                    //       .export
		.coe_f3_out           (a2_f3_out),                                                    //       .export
		.coe_f4_out           (a2_f4_out),                                                    //       .export
		.coe_f5_out           (a2_f5_out),                                                    //       .export
		.coe_f6_out           (a2_f6_out),                                                    //       .export
		.coe_f7_out           (a2_f7_out),                                                    //       .export
		.coe_f_in             (a2_f_in),                                                      //       .export
		.coe_GPIO             (a2_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a3 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a3_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a3_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a3_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a3_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a3_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a3_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a3_f1_oe),                                                     //       .export
		.coe_f2_oe            (a3_f2_oe),                                                     //       .export
		.coe_f3_oe            (a3_f3_oe),                                                     //       .export
		.coe_f4_oe            (a3_f4_oe),                                                     //       .export
		.coe_f5_oe            (a3_f5_oe),                                                     //       .export
		.coe_f6_oe            (a3_f6_oe),                                                     //       .export
		.coe_f7_oe            (a3_f7_oe),                                                     //       .export
		.coe_f0_out           (a3_f0_out),                                                    //       .export
		.coe_f1_out           (a3_f1_out),                                                    //       .export
		.coe_f2_out           (a3_f2_out),                                                    //       .export
		.coe_f3_out           (a3_f3_out),                                                    //       .export
		.coe_f4_out           (a3_f4_out),                                                    //       .export
		.coe_f5_out           (a3_f5_out),                                                    //       .export
		.coe_f6_out           (a3_f6_out),                                                    //       .export
		.coe_f7_out           (a3_f7_out),                                                    //       .export
		.coe_f_in             (a3_f_in),                                                      //       .export
		.coe_GPIO             (a3_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a4 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a4_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a4_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a4_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a4_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a4_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a4_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a4_f1_oe),                                                     //       .export
		.coe_f2_oe            (a4_f2_oe),                                                     //       .export
		.coe_f3_oe            (a4_f3_oe),                                                     //       .export
		.coe_f4_oe            (a4_f4_oe),                                                     //       .export
		.coe_f5_oe            (a4_f5_oe),                                                     //       .export
		.coe_f6_oe            (a4_f6_oe),                                                     //       .export
		.coe_f7_oe            (a4_f7_oe),                                                     //       .export
		.coe_f0_out           (a4_f0_out),                                                    //       .export
		.coe_f1_out           (a4_f1_out),                                                    //       .export
		.coe_f2_out           (a4_f2_out),                                                    //       .export
		.coe_f3_out           (a4_f3_out),                                                    //       .export
		.coe_f4_out           (a4_f4_out),                                                    //       .export
		.coe_f5_out           (a4_f5_out),                                                    //       .export
		.coe_f6_out           (a4_f6_out),                                                    //       .export
		.coe_f7_out           (a4_f7_out),                                                    //       .export
		.coe_f_in             (a4_f_in),                                                      //       .export
		.coe_GPIO             (a4_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a5 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a5_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a5_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a5_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a5_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a5_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a5_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a5_f1_oe),                                                     //       .export
		.coe_f2_oe            (a5_f2_oe),                                                     //       .export
		.coe_f3_oe            (a5_f3_oe),                                                     //       .export
		.coe_f4_oe            (a5_f4_oe),                                                     //       .export
		.coe_f5_oe            (a5_f5_oe),                                                     //       .export
		.coe_f6_oe            (a5_f6_oe),                                                     //       .export
		.coe_f7_oe            (a5_f7_oe),                                                     //       .export
		.coe_f0_out           (a5_f0_out),                                                    //       .export
		.coe_f1_out           (a5_f1_out),                                                    //       .export
		.coe_f2_out           (a5_f2_out),                                                    //       .export
		.coe_f3_out           (a5_f3_out),                                                    //       .export
		.coe_f4_out           (a5_f4_out),                                                    //       .export
		.coe_f5_out           (a5_f5_out),                                                    //       .export
		.coe_f6_out           (a5_f6_out),                                                    //       .export
		.coe_f7_out           (a5_f7_out),                                                    //       .export
		.coe_f_in             (a5_f_in),                                                      //       .export
		.coe_GPIO             (a5_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a6 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a6_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a6_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a6_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a6_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a6_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a6_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a6_f1_oe),                                                     //       .export
		.coe_f2_oe            (a6_f2_oe),                                                     //       .export
		.coe_f3_oe            (a6_f3_oe),                                                     //       .export
		.coe_f4_oe            (a6_f4_oe),                                                     //       .export
		.coe_f5_oe            (a6_f5_oe),                                                     //       .export
		.coe_f6_oe            (a6_f6_oe),                                                     //       .export
		.coe_f7_oe            (a6_f7_oe),                                                     //       .export
		.coe_f0_out           (a6_f0_out),                                                    //       .export
		.coe_f1_out           (a6_f1_out),                                                    //       .export
		.coe_f2_out           (a6_f2_out),                                                    //       .export
		.coe_f3_out           (a6_f3_out),                                                    //       .export
		.coe_f4_out           (a6_f4_out),                                                    //       .export
		.coe_f5_out           (a6_f5_out),                                                    //       .export
		.coe_f6_out           (a6_f6_out),                                                    //       .export
		.coe_f7_out           (a6_f7_out),                                                    //       .export
		.coe_f_in             (a6_f_in),                                                      //       .export
		.coe_GPIO             (a6_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a7 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a7_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a7_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a7_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a7_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a7_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a7_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a7_f1_oe),                                                     //       .export
		.coe_f2_oe            (a7_f2_oe),                                                     //       .export
		.coe_f3_oe            (a7_f3_oe),                                                     //       .export
		.coe_f4_oe            (a7_f4_oe),                                                     //       .export
		.coe_f5_oe            (a7_f5_oe),                                                     //       .export
		.coe_f6_oe            (a7_f6_oe),                                                     //       .export
		.coe_f7_oe            (a7_f7_oe),                                                     //       .export
		.coe_f0_out           (a7_f0_out),                                                    //       .export
		.coe_f1_out           (a7_f1_out),                                                    //       .export
		.coe_f2_out           (a7_f2_out),                                                    //       .export
		.coe_f3_out           (a7_f3_out),                                                    //       .export
		.coe_f4_out           (a7_f4_out),                                                    //       .export
		.coe_f5_out           (a7_f5_out),                                                    //       .export
		.coe_f6_out           (a7_f6_out),                                                    //       .export
		.coe_f7_out           (a7_f7_out),                                                    //       .export
		.coe_f_in             (a7_f_in),                                                      //       .export
		.coe_GPIO             (a7_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a8 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a8_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a8_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a8_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a8_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a8_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a8_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a8_f1_oe),                                                     //       .export
		.coe_f2_oe            (a8_f2_oe),                                                     //       .export
		.coe_f3_oe            (a8_f3_oe),                                                     //       .export
		.coe_f4_oe            (a8_f4_oe),                                                     //       .export
		.coe_f5_oe            (a8_f5_oe),                                                     //       .export
		.coe_f6_oe            (a8_f6_oe),                                                     //       .export
		.coe_f7_oe            (a8_f7_oe),                                                     //       .export
		.coe_f0_out           (a8_f0_out),                                                    //       .export
		.coe_f1_out           (a8_f1_out),                                                    //       .export
		.coe_f2_out           (a8_f2_out),                                                    //       .export
		.coe_f3_out           (a8_f3_out),                                                    //       .export
		.coe_f4_out           (a8_f4_out),                                                    //       .export
		.coe_f5_out           (a8_f5_out),                                                    //       .export
		.coe_f6_out           (a8_f6_out),                                                    //       .export
		.coe_f7_out           (a8_f7_out),                                                    //       .export
		.coe_f_in             (a8_f_in),                                                      //       .export
		.coe_GPIO             (a8_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a9 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a9_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a9_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a9_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a9_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a9_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a9_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a9_f1_oe),                                                     //       .export
		.coe_f2_oe            (a9_f2_oe),                                                     //       .export
		.coe_f3_oe            (a9_f3_oe),                                                     //       .export
		.coe_f4_oe            (a9_f4_oe),                                                     //       .export
		.coe_f5_oe            (a9_f5_oe),                                                     //       .export
		.coe_f6_oe            (a9_f6_oe),                                                     //       .export
		.coe_f7_oe            (a9_f7_oe),                                                     //       .export
		.coe_f0_out           (a9_f0_out),                                                    //       .export
		.coe_f1_out           (a9_f1_out),                                                    //       .export
		.coe_f2_out           (a9_f2_out),                                                    //       .export
		.coe_f3_out           (a9_f3_out),                                                    //       .export
		.coe_f4_out           (a9_f4_out),                                                    //       .export
		.coe_f5_out           (a9_f5_out),                                                    //       .export
		.coe_f6_out           (a9_f6_out),                                                    //       .export
		.coe_f7_out           (a9_f7_out),                                                    //       .export
		.coe_f_in             (a9_f_in),                                                      //       .export
		.coe_GPIO             (a9_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a10 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a10_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a10_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a10_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a10_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a10_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a10_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a10_f1_oe),                                                     //       .export
		.coe_f2_oe            (a10_f2_oe),                                                     //       .export
		.coe_f3_oe            (a10_f3_oe),                                                     //       .export
		.coe_f4_oe            (a10_f4_oe),                                                     //       .export
		.coe_f5_oe            (a10_f5_oe),                                                     //       .export
		.coe_f6_oe            (a10_f6_oe),                                                     //       .export
		.coe_f7_oe            (a10_f7_oe),                                                     //       .export
		.coe_f0_out           (a10_f0_out),                                                    //       .export
		.coe_f1_out           (a10_f1_out),                                                    //       .export
		.coe_f2_out           (a10_f2_out),                                                    //       .export
		.coe_f3_out           (a10_f3_out),                                                    //       .export
		.coe_f4_out           (a10_f4_out),                                                    //       .export
		.coe_f5_out           (a10_f5_out),                                                    //       .export
		.coe_f6_out           (a10_f6_out),                                                    //       .export
		.coe_f7_out           (a10_f7_out),                                                    //       .export
		.coe_f_in             (a10_f_in),                                                      //       .export
		.coe_GPIO             (a10_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a11 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a11_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a11_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a11_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a11_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a11_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a11_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a11_f1_oe),                                                     //       .export
		.coe_f2_oe            (a11_f2_oe),                                                     //       .export
		.coe_f3_oe            (a11_f3_oe),                                                     //       .export
		.coe_f4_oe            (a11_f4_oe),                                                     //       .export
		.coe_f5_oe            (a11_f5_oe),                                                     //       .export
		.coe_f6_oe            (a11_f6_oe),                                                     //       .export
		.coe_f7_oe            (a11_f7_oe),                                                     //       .export
		.coe_f0_out           (a11_f0_out),                                                    //       .export
		.coe_f1_out           (a11_f1_out),                                                    //       .export
		.coe_f2_out           (a11_f2_out),                                                    //       .export
		.coe_f3_out           (a11_f3_out),                                                    //       .export
		.coe_f4_out           (a11_f4_out),                                                    //       .export
		.coe_f5_out           (a11_f5_out),                                                    //       .export
		.coe_f6_out           (a11_f6_out),                                                    //       .export
		.coe_f7_out           (a11_f7_out),                                                    //       .export
		.coe_f_in             (a11_f_in),                                                      //       .export
		.coe_GPIO             (a11_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a12 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a12_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a12_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a12_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a12_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a12_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a12_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a12_f1_oe),                                                     //       .export
		.coe_f2_oe            (a12_f2_oe),                                                     //       .export
		.coe_f3_oe            (a12_f3_oe),                                                     //       .export
		.coe_f4_oe            (a12_f4_oe),                                                     //       .export
		.coe_f5_oe            (a12_f5_oe),                                                     //       .export
		.coe_f6_oe            (a12_f6_oe),                                                     //       .export
		.coe_f7_oe            (a12_f7_oe),                                                     //       .export
		.coe_f0_out           (a12_f0_out),                                                    //       .export
		.coe_f1_out           (a12_f1_out),                                                    //       .export
		.coe_f2_out           (a12_f2_out),                                                    //       .export
		.coe_f3_out           (a12_f3_out),                                                    //       .export
		.coe_f4_out           (a12_f4_out),                                                    //       .export
		.coe_f5_out           (a12_f5_out),                                                    //       .export
		.coe_f6_out           (a12_f6_out),                                                    //       .export
		.coe_f7_out           (a12_f7_out),                                                    //       .export
		.coe_f_in             (a12_f_in),                                                      //       .export
		.coe_GPIO             (a12_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a13 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a13_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a13_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a13_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a13_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a13_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a13_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a13_f1_oe),                                                     //       .export
		.coe_f2_oe            (a13_f2_oe),                                                     //       .export
		.coe_f3_oe            (a13_f3_oe),                                                     //       .export
		.coe_f4_oe            (a13_f4_oe),                                                     //       .export
		.coe_f5_oe            (a13_f5_oe),                                                     //       .export
		.coe_f6_oe            (a13_f6_oe),                                                     //       .export
		.coe_f7_oe            (a13_f7_oe),                                                     //       .export
		.coe_f0_out           (a13_f0_out),                                                    //       .export
		.coe_f1_out           (a13_f1_out),                                                    //       .export
		.coe_f2_out           (a13_f2_out),                                                    //       .export
		.coe_f3_out           (a13_f3_out),                                                    //       .export
		.coe_f4_out           (a13_f4_out),                                                    //       .export
		.coe_f5_out           (a13_f5_out),                                                    //       .export
		.coe_f6_out           (a13_f6_out),                                                    //       .export
		.coe_f7_out           (a13_f7_out),                                                    //       .export
		.coe_f_in             (a13_f_in),                                                      //       .export
		.coe_GPIO             (a13_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a14 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a14_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a14_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a14_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a14_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a14_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a14_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a14_f1_oe),                                                     //       .export
		.coe_f2_oe            (a14_f2_oe),                                                     //       .export
		.coe_f3_oe            (a14_f3_oe),                                                     //       .export
		.coe_f4_oe            (a14_f4_oe),                                                     //       .export
		.coe_f5_oe            (a14_f5_oe),                                                     //       .export
		.coe_f6_oe            (a14_f6_oe),                                                     //       .export
		.coe_f7_oe            (a14_f7_oe),                                                     //       .export
		.coe_f0_out           (a14_f0_out),                                                    //       .export
		.coe_f1_out           (a14_f1_out),                                                    //       .export
		.coe_f2_out           (a14_f2_out),                                                    //       .export
		.coe_f3_out           (a14_f3_out),                                                    //       .export
		.coe_f4_out           (a14_f4_out),                                                    //       .export
		.coe_f5_out           (a14_f5_out),                                                    //       .export
		.coe_f6_out           (a14_f6_out),                                                    //       .export
		.coe_f7_out           (a14_f7_out),                                                    //       .export
		.coe_f_in             (a14_f_in),                                                      //       .export
		.coe_GPIO             (a14_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a15 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a15_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a15_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a15_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a15_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a15_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a15_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a15_f1_oe),                                                     //       .export
		.coe_f2_oe            (a15_f2_oe),                                                     //       .export
		.coe_f3_oe            (a15_f3_oe),                                                     //       .export
		.coe_f4_oe            (a15_f4_oe),                                                     //       .export
		.coe_f5_oe            (a15_f5_oe),                                                     //       .export
		.coe_f6_oe            (a15_f6_oe),                                                     //       .export
		.coe_f7_oe            (a15_f7_oe),                                                     //       .export
		.coe_f0_out           (a15_f0_out),                                                    //       .export
		.coe_f1_out           (a15_f1_out),                                                    //       .export
		.coe_f2_out           (a15_f2_out),                                                    //       .export
		.coe_f3_out           (a15_f3_out),                                                    //       .export
		.coe_f4_out           (a15_f4_out),                                                    //       .export
		.coe_f5_out           (a15_f5_out),                                                    //       .export
		.coe_f6_out           (a15_f6_out),                                                    //       .export
		.coe_f7_out           (a15_f7_out),                                                    //       .export
		.coe_f_in             (a15_f_in),                                                      //       .export
		.coe_GPIO             (a15_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a16 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a16_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a16_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a16_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a16_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a16_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a16_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a16_f1_oe),                                                     //       .export
		.coe_f2_oe            (a16_f2_oe),                                                     //       .export
		.coe_f3_oe            (a16_f3_oe),                                                     //       .export
		.coe_f4_oe            (a16_f4_oe),                                                     //       .export
		.coe_f5_oe            (a16_f5_oe),                                                     //       .export
		.coe_f6_oe            (a16_f6_oe),                                                     //       .export
		.coe_f7_oe            (a16_f7_oe),                                                     //       .export
		.coe_f0_out           (a16_f0_out),                                                    //       .export
		.coe_f1_out           (a16_f1_out),                                                    //       .export
		.coe_f2_out           (a16_f2_out),                                                    //       .export
		.coe_f3_out           (a16_f3_out),                                                    //       .export
		.coe_f4_out           (a16_f4_out),                                                    //       .export
		.coe_f5_out           (a16_f5_out),                                                    //       .export
		.coe_f6_out           (a16_f6_out),                                                    //       .export
		.coe_f7_out           (a16_f7_out),                                                    //       .export
		.coe_f_in             (a16_f_in),                                                      //       .export
		.coe_GPIO             (a16_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a17 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a17_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a17_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a17_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a17_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a17_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a17_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a17_f1_oe),                                                     //       .export
		.coe_f2_oe            (a17_f2_oe),                                                     //       .export
		.coe_f3_oe            (a17_f3_oe),                                                     //       .export
		.coe_f4_oe            (a17_f4_oe),                                                     //       .export
		.coe_f5_oe            (a17_f5_oe),                                                     //       .export
		.coe_f6_oe            (a17_f6_oe),                                                     //       .export
		.coe_f7_oe            (a17_f7_oe),                                                     //       .export
		.coe_f0_out           (a17_f0_out),                                                    //       .export
		.coe_f1_out           (a17_f1_out),                                                    //       .export
		.coe_f2_out           (a17_f2_out),                                                    //       .export
		.coe_f3_out           (a17_f3_out),                                                    //       .export
		.coe_f4_out           (a17_f4_out),                                                    //       .export
		.coe_f5_out           (a17_f5_out),                                                    //       .export
		.coe_f6_out           (a17_f6_out),                                                    //       .export
		.coe_f7_out           (a17_f7_out),                                                    //       .export
		.coe_f_in             (a17_f_in),                                                      //       .export
		.coe_GPIO             (a17_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a18 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a18_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a18_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a18_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a18_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a18_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a18_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a18_f1_oe),                                                     //       .export
		.coe_f2_oe            (a18_f2_oe),                                                     //       .export
		.coe_f3_oe            (a18_f3_oe),                                                     //       .export
		.coe_f4_oe            (a18_f4_oe),                                                     //       .export
		.coe_f5_oe            (a18_f5_oe),                                                     //       .export
		.coe_f6_oe            (a18_f6_oe),                                                     //       .export
		.coe_f7_oe            (a18_f7_oe),                                                     //       .export
		.coe_f0_out           (a18_f0_out),                                                    //       .export
		.coe_f1_out           (a18_f1_out),                                                    //       .export
		.coe_f2_out           (a18_f2_out),                                                    //       .export
		.coe_f3_out           (a18_f3_out),                                                    //       .export
		.coe_f4_out           (a18_f4_out),                                                    //       .export
		.coe_f5_out           (a18_f5_out),                                                    //       .export
		.coe_f6_out           (a18_f6_out),                                                    //       .export
		.coe_f7_out           (a18_f7_out),                                                    //       .export
		.coe_f_in             (a18_f_in),                                                      //       .export
		.coe_GPIO             (a18_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a19 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a19_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a19_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a19_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a19_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a19_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a19_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a19_f1_oe),                                                     //       .export
		.coe_f2_oe            (a19_f2_oe),                                                     //       .export
		.coe_f3_oe            (a19_f3_oe),                                                     //       .export
		.coe_f4_oe            (a19_f4_oe),                                                     //       .export
		.coe_f5_oe            (a19_f5_oe),                                                     //       .export
		.coe_f6_oe            (a19_f6_oe),                                                     //       .export
		.coe_f7_oe            (a19_f7_oe),                                                     //       .export
		.coe_f0_out           (a19_f0_out),                                                    //       .export
		.coe_f1_out           (a19_f1_out),                                                    //       .export
		.coe_f2_out           (a19_f2_out),                                                    //       .export
		.coe_f3_out           (a19_f3_out),                                                    //       .export
		.coe_f4_out           (a19_f4_out),                                                    //       .export
		.coe_f5_out           (a19_f5_out),                                                    //       .export
		.coe_f6_out           (a19_f6_out),                                                    //       .export
		.coe_f7_out           (a19_f7_out),                                                    //       .export
		.coe_f_in             (a19_f_in),                                                      //       .export
		.coe_GPIO             (a19_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a20 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a20_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a20_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a20_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a20_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a20_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a20_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a20_f1_oe),                                                     //       .export
		.coe_f2_oe            (a20_f2_oe),                                                     //       .export
		.coe_f3_oe            (a20_f3_oe),                                                     //       .export
		.coe_f4_oe            (a20_f4_oe),                                                     //       .export
		.coe_f5_oe            (a20_f5_oe),                                                     //       .export
		.coe_f6_oe            (a20_f6_oe),                                                     //       .export
		.coe_f7_oe            (a20_f7_oe),                                                     //       .export
		.coe_f0_out           (a20_f0_out),                                                    //       .export
		.coe_f1_out           (a20_f1_out),                                                    //       .export
		.coe_f2_out           (a20_f2_out),                                                    //       .export
		.coe_f3_out           (a20_f3_out),                                                    //       .export
		.coe_f4_out           (a20_f4_out),                                                    //       .export
		.coe_f5_out           (a20_f5_out),                                                    //       .export
		.coe_f6_out           (a20_f6_out),                                                    //       .export
		.coe_f7_out           (a20_f7_out),                                                    //       .export
		.coe_f_in             (a20_f_in),                                                      //       .export
		.coe_GPIO             (a20_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a21 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a21_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a21_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a21_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a21_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a21_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a21_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a21_f1_oe),                                                     //       .export
		.coe_f2_oe            (a21_f2_oe),                                                     //       .export
		.coe_f3_oe            (a21_f3_oe),                                                     //       .export
		.coe_f4_oe            (a21_f4_oe),                                                     //       .export
		.coe_f5_oe            (a21_f5_oe),                                                     //       .export
		.coe_f6_oe            (a21_f6_oe),                                                     //       .export
		.coe_f7_oe            (a21_f7_oe),                                                     //       .export
		.coe_f0_out           (a21_f0_out),                                                    //       .export
		.coe_f1_out           (a21_f1_out),                                                    //       .export
		.coe_f2_out           (a21_f2_out),                                                    //       .export
		.coe_f3_out           (a21_f3_out),                                                    //       .export
		.coe_f4_out           (a21_f4_out),                                                    //       .export
		.coe_f5_out           (a21_f5_out),                                                    //       .export
		.coe_f6_out           (a21_f6_out),                                                    //       .export
		.coe_f7_out           (a21_f7_out),                                                    //       .export
		.coe_f_in             (a21_f_in),                                                      //       .export
		.coe_GPIO             (a21_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a22 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a22_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a22_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a22_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a22_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a22_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a22_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a22_f1_oe),                                                     //       .export
		.coe_f2_oe            (a22_f2_oe),                                                     //       .export
		.coe_f3_oe            (a22_f3_oe),                                                     //       .export
		.coe_f4_oe            (a22_f4_oe),                                                     //       .export
		.coe_f5_oe            (a22_f5_oe),                                                     //       .export
		.coe_f6_oe            (a22_f6_oe),                                                     //       .export
		.coe_f7_oe            (a22_f7_oe),                                                     //       .export
		.coe_f0_out           (a22_f0_out),                                                    //       .export
		.coe_f1_out           (a22_f1_out),                                                    //       .export
		.coe_f2_out           (a22_f2_out),                                                    //       .export
		.coe_f3_out           (a22_f3_out),                                                    //       .export
		.coe_f4_out           (a22_f4_out),                                                    //       .export
		.coe_f5_out           (a22_f5_out),                                                    //       .export
		.coe_f6_out           (a22_f6_out),                                                    //       .export
		.coe_f7_out           (a22_f7_out),                                                    //       .export
		.coe_f_in             (a22_f_in),                                                      //       .export
		.coe_GPIO             (a22_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a23 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a23_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a23_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a23_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a23_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a23_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a23_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a23_f1_oe),                                                     //       .export
		.coe_f2_oe            (a23_f2_oe),                                                     //       .export
		.coe_f3_oe            (a23_f3_oe),                                                     //       .export
		.coe_f4_oe            (a23_f4_oe),                                                     //       .export
		.coe_f5_oe            (a23_f5_oe),                                                     //       .export
		.coe_f6_oe            (a23_f6_oe),                                                     //       .export
		.coe_f7_oe            (a23_f7_oe),                                                     //       .export
		.coe_f0_out           (a23_f0_out),                                                    //       .export
		.coe_f1_out           (a23_f1_out),                                                    //       .export
		.coe_f2_out           (a23_f2_out),                                                    //       .export
		.coe_f3_out           (a23_f3_out),                                                    //       .export
		.coe_f4_out           (a23_f4_out),                                                    //       .export
		.coe_f5_out           (a23_f5_out),                                                    //       .export
		.coe_f6_out           (a23_f6_out),                                                    //       .export
		.coe_f7_out           (a23_f7_out),                                                    //       .export
		.coe_f_in             (a23_f_in),                                                      //       .export
		.coe_GPIO             (a23_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a24 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a24_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a24_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a24_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a24_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a24_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a24_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a24_f1_oe),                                                     //       .export
		.coe_f2_oe            (a24_f2_oe),                                                     //       .export
		.coe_f3_oe            (a24_f3_oe),                                                     //       .export
		.coe_f4_oe            (a24_f4_oe),                                                     //       .export
		.coe_f5_oe            (a24_f5_oe),                                                     //       .export
		.coe_f6_oe            (a24_f6_oe),                                                     //       .export
		.coe_f7_oe            (a24_f7_oe),                                                     //       .export
		.coe_f0_out           (a24_f0_out),                                                    //       .export
		.coe_f1_out           (a24_f1_out),                                                    //       .export
		.coe_f2_out           (a24_f2_out),                                                    //       .export
		.coe_f3_out           (a24_f3_out),                                                    //       .export
		.coe_f4_out           (a24_f4_out),                                                    //       .export
		.coe_f5_out           (a24_f5_out),                                                    //       .export
		.coe_f6_out           (a24_f6_out),                                                    //       .export
		.coe_f7_out           (a24_f7_out),                                                    //       .export
		.coe_f_in             (a24_f_in),                                                      //       .export
		.coe_GPIO             (a24_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_a25 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_a25_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_a25_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_a25_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_a25_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_a25_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (a25_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (a25_f1_oe),                                                     //       .export
		.coe_f2_oe            (a25_f2_oe),                                                     //       .export
		.coe_f3_oe            (a25_f3_oe),                                                     //       .export
		.coe_f4_oe            (a25_f4_oe),                                                     //       .export
		.coe_f5_oe            (a25_f5_oe),                                                     //       .export
		.coe_f6_oe            (a25_f6_oe),                                                     //       .export
		.coe_f7_oe            (a25_f7_oe),                                                     //       .export
		.coe_f0_out           (a25_f0_out),                                                    //       .export
		.coe_f1_out           (a25_f1_out),                                                    //       .export
		.coe_f2_out           (a25_f2_out),                                                    //       .export
		.coe_f3_out           (a25_f3_out),                                                    //       .export
		.coe_f4_out           (a25_f4_out),                                                    //       .export
		.coe_f5_out           (a25_f5_out),                                                    //       .export
		.coe_f6_out           (a25_f6_out),                                                    //       .export
		.coe_f7_out           (a25_f7_out),                                                    //       .export
		.coe_f_in             (a25_f_in),                                                      //       .export
		.coe_GPIO             (a25_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b0 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b0_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b0_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b0_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b0_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b0_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b0_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b0_f1_oe),                                                     //       .export
		.coe_f2_oe            (b0_f2_oe),                                                     //       .export
		.coe_f3_oe            (b0_f3_oe),                                                     //       .export
		.coe_f4_oe            (b0_f4_oe),                                                     //       .export
		.coe_f5_oe            (b0_f5_oe),                                                     //       .export
		.coe_f6_oe            (b0_f6_oe),                                                     //       .export
		.coe_f7_oe            (b0_f7_oe),                                                     //       .export
		.coe_f0_out           (b0_f0_out),                                                    //       .export
		.coe_f1_out           (b0_f1_out),                                                    //       .export
		.coe_f2_out           (b0_f2_out),                                                    //       .export
		.coe_f3_out           (b0_f3_out),                                                    //       .export
		.coe_f4_out           (b0_f4_out),                                                    //       .export
		.coe_f5_out           (b0_f5_out),                                                    //       .export
		.coe_f6_out           (b0_f6_out),                                                    //       .export
		.coe_f7_out           (b0_f7_out),                                                    //       .export
		.coe_f_in             (b0_f_in),                                                      //       .export
		.coe_GPIO             (b0_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b1 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b1_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b1_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b1_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b1_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b1_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b1_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b1_f1_oe),                                                     //       .export
		.coe_f2_oe            (b1_f2_oe),                                                     //       .export
		.coe_f3_oe            (b1_f3_oe),                                                     //       .export
		.coe_f4_oe            (b1_f4_oe),                                                     //       .export
		.coe_f5_oe            (b1_f5_oe),                                                     //       .export
		.coe_f6_oe            (b1_f6_oe),                                                     //       .export
		.coe_f7_oe            (b1_f7_oe),                                                     //       .export
		.coe_f0_out           (b1_f0_out),                                                    //       .export
		.coe_f1_out           (b1_f1_out),                                                    //       .export
		.coe_f2_out           (b1_f2_out),                                                    //       .export
		.coe_f3_out           (b1_f3_out),                                                    //       .export
		.coe_f4_out           (b1_f4_out),                                                    //       .export
		.coe_f5_out           (b1_f5_out),                                                    //       .export
		.coe_f6_out           (b1_f6_out),                                                    //       .export
		.coe_f7_out           (b1_f7_out),                                                    //       .export
		.coe_f_in             (b1_f_in),                                                      //       .export
		.coe_GPIO             (b1_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b2 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b2_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b2_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b2_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b2_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b2_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b2_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b2_f1_oe),                                                     //       .export
		.coe_f2_oe            (b2_f2_oe),                                                     //       .export
		.coe_f3_oe            (b2_f3_oe),                                                     //       .export
		.coe_f4_oe            (b2_f4_oe),                                                     //       .export
		.coe_f5_oe            (b2_f5_oe),                                                     //       .export
		.coe_f6_oe            (b2_f6_oe),                                                     //       .export
		.coe_f7_oe            (b2_f7_oe),                                                     //       .export
		.coe_f0_out           (b2_f0_out),                                                    //       .export
		.coe_f1_out           (b2_f1_out),                                                    //       .export
		.coe_f2_out           (b2_f2_out),                                                    //       .export
		.coe_f3_out           (b2_f3_out),                                                    //       .export
		.coe_f4_out           (b2_f4_out),                                                    //       .export
		.coe_f5_out           (b2_f5_out),                                                    //       .export
		.coe_f6_out           (b2_f6_out),                                                    //       .export
		.coe_f7_out           (b2_f7_out),                                                    //       .export
		.coe_f_in             (b2_f_in),                                                      //       .export
		.coe_GPIO             (b2_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b3 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b3_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b3_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b3_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b3_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b3_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b3_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b3_f1_oe),                                                     //       .export
		.coe_f2_oe            (b3_f2_oe),                                                     //       .export
		.coe_f3_oe            (b3_f3_oe),                                                     //       .export
		.coe_f4_oe            (b3_f4_oe),                                                     //       .export
		.coe_f5_oe            (b3_f5_oe),                                                     //       .export
		.coe_f6_oe            (b3_f6_oe),                                                     //       .export
		.coe_f7_oe            (b3_f7_oe),                                                     //       .export
		.coe_f0_out           (b3_f0_out),                                                    //       .export
		.coe_f1_out           (b3_f1_out),                                                    //       .export
		.coe_f2_out           (b3_f2_out),                                                    //       .export
		.coe_f3_out           (b3_f3_out),                                                    //       .export
		.coe_f4_out           (b3_f4_out),                                                    //       .export
		.coe_f5_out           (b3_f5_out),                                                    //       .export
		.coe_f6_out           (b3_f6_out),                                                    //       .export
		.coe_f7_out           (b3_f7_out),                                                    //       .export
		.coe_f_in             (b3_f_in),                                                      //       .export
		.coe_GPIO             (b3_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b4 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b4_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b4_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b4_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b4_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b4_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b4_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b4_f1_oe),                                                     //       .export
		.coe_f2_oe            (b4_f2_oe),                                                     //       .export
		.coe_f3_oe            (b4_f3_oe),                                                     //       .export
		.coe_f4_oe            (b4_f4_oe),                                                     //       .export
		.coe_f5_oe            (b4_f5_oe),                                                     //       .export
		.coe_f6_oe            (b4_f6_oe),                                                     //       .export
		.coe_f7_oe            (b4_f7_oe),                                                     //       .export
		.coe_f0_out           (b4_f0_out),                                                    //       .export
		.coe_f1_out           (b4_f1_out),                                                    //       .export
		.coe_f2_out           (b4_f2_out),                                                    //       .export
		.coe_f3_out           (b4_f3_out),                                                    //       .export
		.coe_f4_out           (b4_f4_out),                                                    //       .export
		.coe_f5_out           (b4_f5_out),                                                    //       .export
		.coe_f6_out           (b4_f6_out),                                                    //       .export
		.coe_f7_out           (b4_f7_out),                                                    //       .export
		.coe_f_in             (b4_f_in),                                                      //       .export
		.coe_GPIO             (b4_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b5 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b5_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b5_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b5_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b5_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b5_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b5_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b5_f1_oe),                                                     //       .export
		.coe_f2_oe            (b5_f2_oe),                                                     //       .export
		.coe_f3_oe            (b5_f3_oe),                                                     //       .export
		.coe_f4_oe            (b5_f4_oe),                                                     //       .export
		.coe_f5_oe            (b5_f5_oe),                                                     //       .export
		.coe_f6_oe            (b5_f6_oe),                                                     //       .export
		.coe_f7_oe            (b5_f7_oe),                                                     //       .export
		.coe_f0_out           (b5_f0_out),                                                    //       .export
		.coe_f1_out           (b5_f1_out),                                                    //       .export
		.coe_f2_out           (b5_f2_out),                                                    //       .export
		.coe_f3_out           (b5_f3_out),                                                    //       .export
		.coe_f4_out           (b5_f4_out),                                                    //       .export
		.coe_f5_out           (b5_f5_out),                                                    //       .export
		.coe_f6_out           (b5_f6_out),                                                    //       .export
		.coe_f7_out           (b5_f7_out),                                                    //       .export
		.coe_f_in             (b5_f_in),                                                      //       .export
		.coe_GPIO             (b5_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b6 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b6_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b6_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b6_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b6_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b6_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b6_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b6_f1_oe),                                                     //       .export
		.coe_f2_oe            (b6_f2_oe),                                                     //       .export
		.coe_f3_oe            (b6_f3_oe),                                                     //       .export
		.coe_f4_oe            (b6_f4_oe),                                                     //       .export
		.coe_f5_oe            (b6_f5_oe),                                                     //       .export
		.coe_f6_oe            (b6_f6_oe),                                                     //       .export
		.coe_f7_oe            (b6_f7_oe),                                                     //       .export
		.coe_f0_out           (b6_f0_out),                                                    //       .export
		.coe_f1_out           (b6_f1_out),                                                    //       .export
		.coe_f2_out           (b6_f2_out),                                                    //       .export
		.coe_f3_out           (b6_f3_out),                                                    //       .export
		.coe_f4_out           (b6_f4_out),                                                    //       .export
		.coe_f5_out           (b6_f5_out),                                                    //       .export
		.coe_f6_out           (b6_f6_out),                                                    //       .export
		.coe_f7_out           (b6_f7_out),                                                    //       .export
		.coe_f_in             (b6_f_in),                                                      //       .export
		.coe_GPIO             (b6_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b7 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b7_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b7_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b7_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b7_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b7_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b7_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b7_f1_oe),                                                     //       .export
		.coe_f2_oe            (b7_f2_oe),                                                     //       .export
		.coe_f3_oe            (b7_f3_oe),                                                     //       .export
		.coe_f4_oe            (b7_f4_oe),                                                     //       .export
		.coe_f5_oe            (b7_f5_oe),                                                     //       .export
		.coe_f6_oe            (b7_f6_oe),                                                     //       .export
		.coe_f7_oe            (b7_f7_oe),                                                     //       .export
		.coe_f0_out           (b7_f0_out),                                                    //       .export
		.coe_f1_out           (b7_f1_out),                                                    //       .export
		.coe_f2_out           (b7_f2_out),                                                    //       .export
		.coe_f3_out           (b7_f3_out),                                                    //       .export
		.coe_f4_out           (b7_f4_out),                                                    //       .export
		.coe_f5_out           (b7_f5_out),                                                    //       .export
		.coe_f6_out           (b7_f6_out),                                                    //       .export
		.coe_f7_out           (b7_f7_out),                                                    //       .export
		.coe_f_in             (b7_f_in),                                                      //       .export
		.coe_GPIO             (b7_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b8 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b8_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b8_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b8_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b8_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b8_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b8_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b8_f1_oe),                                                     //       .export
		.coe_f2_oe            (b8_f2_oe),                                                     //       .export
		.coe_f3_oe            (b8_f3_oe),                                                     //       .export
		.coe_f4_oe            (b8_f4_oe),                                                     //       .export
		.coe_f5_oe            (b8_f5_oe),                                                     //       .export
		.coe_f6_oe            (b8_f6_oe),                                                     //       .export
		.coe_f7_oe            (b8_f7_oe),                                                     //       .export
		.coe_f0_out           (b8_f0_out),                                                    //       .export
		.coe_f1_out           (b8_f1_out),                                                    //       .export
		.coe_f2_out           (b8_f2_out),                                                    //       .export
		.coe_f3_out           (b8_f3_out),                                                    //       .export
		.coe_f4_out           (b8_f4_out),                                                    //       .export
		.coe_f5_out           (b8_f5_out),                                                    //       .export
		.coe_f6_out           (b8_f6_out),                                                    //       .export
		.coe_f7_out           (b8_f7_out),                                                    //       .export
		.coe_f_in             (b8_f_in),                                                      //       .export
		.coe_GPIO             (b8_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b9 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b9_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b9_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b9_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b9_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b9_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b9_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b9_f1_oe),                                                     //       .export
		.coe_f2_oe            (b9_f2_oe),                                                     //       .export
		.coe_f3_oe            (b9_f3_oe),                                                     //       .export
		.coe_f4_oe            (b9_f4_oe),                                                     //       .export
		.coe_f5_oe            (b9_f5_oe),                                                     //       .export
		.coe_f6_oe            (b9_f6_oe),                                                     //       .export
		.coe_f7_oe            (b9_f7_oe),                                                     //       .export
		.coe_f0_out           (b9_f0_out),                                                    //       .export
		.coe_f1_out           (b9_f1_out),                                                    //       .export
		.coe_f2_out           (b9_f2_out),                                                    //       .export
		.coe_f3_out           (b9_f3_out),                                                    //       .export
		.coe_f4_out           (b9_f4_out),                                                    //       .export
		.coe_f5_out           (b9_f5_out),                                                    //       .export
		.coe_f6_out           (b9_f6_out),                                                    //       .export
		.coe_f7_out           (b9_f7_out),                                                    //       .export
		.coe_f_in             (b9_f_in),                                                      //       .export
		.coe_GPIO             (b9_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b10 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b10_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b10_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b10_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b10_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b10_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b10_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b10_f1_oe),                                                     //       .export
		.coe_f2_oe            (b10_f2_oe),                                                     //       .export
		.coe_f3_oe            (b10_f3_oe),                                                     //       .export
		.coe_f4_oe            (b10_f4_oe),                                                     //       .export
		.coe_f5_oe            (b10_f5_oe),                                                     //       .export
		.coe_f6_oe            (b10_f6_oe),                                                     //       .export
		.coe_f7_oe            (b10_f7_oe),                                                     //       .export
		.coe_f0_out           (b10_f0_out),                                                    //       .export
		.coe_f1_out           (b10_f1_out),                                                    //       .export
		.coe_f2_out           (b10_f2_out),                                                    //       .export
		.coe_f3_out           (b10_f3_out),                                                    //       .export
		.coe_f4_out           (b10_f4_out),                                                    //       .export
		.coe_f5_out           (b10_f5_out),                                                    //       .export
		.coe_f6_out           (b10_f6_out),                                                    //       .export
		.coe_f7_out           (b10_f7_out),                                                    //       .export
		.coe_f_in             (b10_f_in),                                                      //       .export
		.coe_GPIO             (b10_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b11 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b11_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b11_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b11_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b11_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b11_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b11_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b11_f1_oe),                                                     //       .export
		.coe_f2_oe            (b11_f2_oe),                                                     //       .export
		.coe_f3_oe            (b11_f3_oe),                                                     //       .export
		.coe_f4_oe            (b11_f4_oe),                                                     //       .export
		.coe_f5_oe            (b11_f5_oe),                                                     //       .export
		.coe_f6_oe            (b11_f6_oe),                                                     //       .export
		.coe_f7_oe            (b11_f7_oe),                                                     //       .export
		.coe_f0_out           (b11_f0_out),                                                    //       .export
		.coe_f1_out           (b11_f1_out),                                                    //       .export
		.coe_f2_out           (b11_f2_out),                                                    //       .export
		.coe_f3_out           (b11_f3_out),                                                    //       .export
		.coe_f4_out           (b11_f4_out),                                                    //       .export
		.coe_f5_out           (b11_f5_out),                                                    //       .export
		.coe_f6_out           (b11_f6_out),                                                    //       .export
		.coe_f7_out           (b11_f7_out),                                                    //       .export
		.coe_f_in             (b11_f_in),                                                      //       .export
		.coe_GPIO             (b11_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b12 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b12_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b12_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b12_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b12_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b12_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b12_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b12_f1_oe),                                                     //       .export
		.coe_f2_oe            (b12_f2_oe),                                                     //       .export
		.coe_f3_oe            (b12_f3_oe),                                                     //       .export
		.coe_f4_oe            (b12_f4_oe),                                                     //       .export
		.coe_f5_oe            (b12_f5_oe),                                                     //       .export
		.coe_f6_oe            (b12_f6_oe),                                                     //       .export
		.coe_f7_oe            (b12_f7_oe),                                                     //       .export
		.coe_f0_out           (b12_f0_out),                                                    //       .export
		.coe_f1_out           (b12_f1_out),                                                    //       .export
		.coe_f2_out           (b12_f2_out),                                                    //       .export
		.coe_f3_out           (b12_f3_out),                                                    //       .export
		.coe_f4_out           (b12_f4_out),                                                    //       .export
		.coe_f5_out           (b12_f5_out),                                                    //       .export
		.coe_f6_out           (b12_f6_out),                                                    //       .export
		.coe_f7_out           (b12_f7_out),                                                    //       .export
		.coe_f_in             (b12_f_in),                                                      //       .export
		.coe_GPIO             (b12_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b13 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b13_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b13_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b13_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b13_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b13_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b13_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b13_f1_oe),                                                     //       .export
		.coe_f2_oe            (b13_f2_oe),                                                     //       .export
		.coe_f3_oe            (b13_f3_oe),                                                     //       .export
		.coe_f4_oe            (b13_f4_oe),                                                     //       .export
		.coe_f5_oe            (b13_f5_oe),                                                     //       .export
		.coe_f6_oe            (b13_f6_oe),                                                     //       .export
		.coe_f7_oe            (b13_f7_oe),                                                     //       .export
		.coe_f0_out           (b13_f0_out),                                                    //       .export
		.coe_f1_out           (b13_f1_out),                                                    //       .export
		.coe_f2_out           (b13_f2_out),                                                    //       .export
		.coe_f3_out           (b13_f3_out),                                                    //       .export
		.coe_f4_out           (b13_f4_out),                                                    //       .export
		.coe_f5_out           (b13_f5_out),                                                    //       .export
		.coe_f6_out           (b13_f6_out),                                                    //       .export
		.coe_f7_out           (b13_f7_out),                                                    //       .export
		.coe_f_in             (b13_f_in),                                                      //       .export
		.coe_GPIO             (b13_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b14 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b14_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b14_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b14_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b14_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b14_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b14_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b14_f1_oe),                                                     //       .export
		.coe_f2_oe            (b14_f2_oe),                                                     //       .export
		.coe_f3_oe            (b14_f3_oe),                                                     //       .export
		.coe_f4_oe            (b14_f4_oe),                                                     //       .export
		.coe_f5_oe            (b14_f5_oe),                                                     //       .export
		.coe_f6_oe            (b14_f6_oe),                                                     //       .export
		.coe_f7_oe            (b14_f7_oe),                                                     //       .export
		.coe_f0_out           (b14_f0_out),                                                    //       .export
		.coe_f1_out           (b14_f1_out),                                                    //       .export
		.coe_f2_out           (b14_f2_out),                                                    //       .export
		.coe_f3_out           (b14_f3_out),                                                    //       .export
		.coe_f4_out           (b14_f4_out),                                                    //       .export
		.coe_f5_out           (b14_f5_out),                                                    //       .export
		.coe_f6_out           (b14_f6_out),                                                    //       .export
		.coe_f7_out           (b14_f7_out),                                                    //       .export
		.coe_f_in             (b14_f_in),                                                      //       .export
		.coe_GPIO             (b14_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b15 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b15_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b15_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b15_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b15_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b15_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b15_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b15_f1_oe),                                                     //       .export
		.coe_f2_oe            (b15_f2_oe),                                                     //       .export
		.coe_f3_oe            (b15_f3_oe),                                                     //       .export
		.coe_f4_oe            (b15_f4_oe),                                                     //       .export
		.coe_f5_oe            (b15_f5_oe),                                                     //       .export
		.coe_f6_oe            (b15_f6_oe),                                                     //       .export
		.coe_f7_oe            (b15_f7_oe),                                                     //       .export
		.coe_f0_out           (b15_f0_out),                                                    //       .export
		.coe_f1_out           (b15_f1_out),                                                    //       .export
		.coe_f2_out           (b15_f2_out),                                                    //       .export
		.coe_f3_out           (b15_f3_out),                                                    //       .export
		.coe_f4_out           (b15_f4_out),                                                    //       .export
		.coe_f5_out           (b15_f5_out),                                                    //       .export
		.coe_f6_out           (b15_f6_out),                                                    //       .export
		.coe_f7_out           (b15_f7_out),                                                    //       .export
		.coe_f_in             (b15_f_in),                                                      //       .export
		.coe_GPIO             (b15_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b16 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b16_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b16_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b16_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b16_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b16_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b16_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b16_f1_oe),                                                     //       .export
		.coe_f2_oe            (b16_f2_oe),                                                     //       .export
		.coe_f3_oe            (b16_f3_oe),                                                     //       .export
		.coe_f4_oe            (b16_f4_oe),                                                     //       .export
		.coe_f5_oe            (b16_f5_oe),                                                     //       .export
		.coe_f6_oe            (b16_f6_oe),                                                     //       .export
		.coe_f7_oe            (b16_f7_oe),                                                     //       .export
		.coe_f0_out           (b16_f0_out),                                                    //       .export
		.coe_f1_out           (b16_f1_out),                                                    //       .export
		.coe_f2_out           (b16_f2_out),                                                    //       .export
		.coe_f3_out           (b16_f3_out),                                                    //       .export
		.coe_f4_out           (b16_f4_out),                                                    //       .export
		.coe_f5_out           (b16_f5_out),                                                    //       .export
		.coe_f6_out           (b16_f6_out),                                                    //       .export
		.coe_f7_out           (b16_f7_out),                                                    //       .export
		.coe_f_in             (b16_f_in),                                                      //       .export
		.coe_GPIO             (b16_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b17 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b17_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b17_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b17_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b17_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b17_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b17_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b17_f1_oe),                                                     //       .export
		.coe_f2_oe            (b17_f2_oe),                                                     //       .export
		.coe_f3_oe            (b17_f3_oe),                                                     //       .export
		.coe_f4_oe            (b17_f4_oe),                                                     //       .export
		.coe_f5_oe            (b17_f5_oe),                                                     //       .export
		.coe_f6_oe            (b17_f6_oe),                                                     //       .export
		.coe_f7_oe            (b17_f7_oe),                                                     //       .export
		.coe_f0_out           (b17_f0_out),                                                    //       .export
		.coe_f1_out           (b17_f1_out),                                                    //       .export
		.coe_f2_out           (b17_f2_out),                                                    //       .export
		.coe_f3_out           (b17_f3_out),                                                    //       .export
		.coe_f4_out           (b17_f4_out),                                                    //       .export
		.coe_f5_out           (b17_f5_out),                                                    //       .export
		.coe_f6_out           (b17_f6_out),                                                    //       .export
		.coe_f7_out           (b17_f7_out),                                                    //       .export
		.coe_f_in             (b17_f_in),                                                      //       .export
		.coe_GPIO             (b17_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b18 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b18_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b18_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b18_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b18_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b18_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b18_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b18_f1_oe),                                                     //       .export
		.coe_f2_oe            (b18_f2_oe),                                                     //       .export
		.coe_f3_oe            (b18_f3_oe),                                                     //       .export
		.coe_f4_oe            (b18_f4_oe),                                                     //       .export
		.coe_f5_oe            (b18_f5_oe),                                                     //       .export
		.coe_f6_oe            (b18_f6_oe),                                                     //       .export
		.coe_f7_oe            (b18_f7_oe),                                                     //       .export
		.coe_f0_out           (b18_f0_out),                                                    //       .export
		.coe_f1_out           (b18_f1_out),                                                    //       .export
		.coe_f2_out           (b18_f2_out),                                                    //       .export
		.coe_f3_out           (b18_f3_out),                                                    //       .export
		.coe_f4_out           (b18_f4_out),                                                    //       .export
		.coe_f5_out           (b18_f5_out),                                                    //       .export
		.coe_f6_out           (b18_f6_out),                                                    //       .export
		.coe_f7_out           (b18_f7_out),                                                    //       .export
		.coe_f_in             (b18_f_in),                                                      //       .export
		.coe_GPIO             (b18_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b19 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b19_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b19_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b19_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b19_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b19_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b19_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b19_f1_oe),                                                     //       .export
		.coe_f2_oe            (b19_f2_oe),                                                     //       .export
		.coe_f3_oe            (b19_f3_oe),                                                     //       .export
		.coe_f4_oe            (b19_f4_oe),                                                     //       .export
		.coe_f5_oe            (b19_f5_oe),                                                     //       .export
		.coe_f6_oe            (b19_f6_oe),                                                     //       .export
		.coe_f7_oe            (b19_f7_oe),                                                     //       .export
		.coe_f0_out           (b19_f0_out),                                                    //       .export
		.coe_f1_out           (b19_f1_out),                                                    //       .export
		.coe_f2_out           (b19_f2_out),                                                    //       .export
		.coe_f3_out           (b19_f3_out),                                                    //       .export
		.coe_f4_out           (b19_f4_out),                                                    //       .export
		.coe_f5_out           (b19_f5_out),                                                    //       .export
		.coe_f6_out           (b19_f6_out),                                                    //       .export
		.coe_f7_out           (b19_f7_out),                                                    //       .export
		.coe_f_in             (b19_f_in),                                                      //       .export
		.coe_GPIO             (b19_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b20 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b20_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b20_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b20_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b20_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b20_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b20_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b20_f1_oe),                                                     //       .export
		.coe_f2_oe            (b20_f2_oe),                                                     //       .export
		.coe_f3_oe            (b20_f3_oe),                                                     //       .export
		.coe_f4_oe            (b20_f4_oe),                                                     //       .export
		.coe_f5_oe            (b20_f5_oe),                                                     //       .export
		.coe_f6_oe            (b20_f6_oe),                                                     //       .export
		.coe_f7_oe            (b20_f7_oe),                                                     //       .export
		.coe_f0_out           (b20_f0_out),                                                    //       .export
		.coe_f1_out           (b20_f1_out),                                                    //       .export
		.coe_f2_out           (b20_f2_out),                                                    //       .export
		.coe_f3_out           (b20_f3_out),                                                    //       .export
		.coe_f4_out           (b20_f4_out),                                                    //       .export
		.coe_f5_out           (b20_f5_out),                                                    //       .export
		.coe_f6_out           (b20_f6_out),                                                    //       .export
		.coe_f7_out           (b20_f7_out),                                                    //       .export
		.coe_f_in             (b20_f_in),                                                      //       .export
		.coe_GPIO             (b20_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b21 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b21_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b21_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b21_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b21_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b21_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b21_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b21_f1_oe),                                                     //       .export
		.coe_f2_oe            (b21_f2_oe),                                                     //       .export
		.coe_f3_oe            (b21_f3_oe),                                                     //       .export
		.coe_f4_oe            (b21_f4_oe),                                                     //       .export
		.coe_f5_oe            (b21_f5_oe),                                                     //       .export
		.coe_f6_oe            (b21_f6_oe),                                                     //       .export
		.coe_f7_oe            (b21_f7_oe),                                                     //       .export
		.coe_f0_out           (b21_f0_out),                                                    //       .export
		.coe_f1_out           (b21_f1_out),                                                    //       .export
		.coe_f2_out           (b21_f2_out),                                                    //       .export
		.coe_f3_out           (b21_f3_out),                                                    //       .export
		.coe_f4_out           (b21_f4_out),                                                    //       .export
		.coe_f5_out           (b21_f5_out),                                                    //       .export
		.coe_f6_out           (b21_f6_out),                                                    //       .export
		.coe_f7_out           (b21_f7_out),                                                    //       .export
		.coe_f_in             (b21_f_in),                                                      //       .export
		.coe_GPIO             (b21_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b22 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b22_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b22_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b22_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b22_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b22_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b22_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b22_f1_oe),                                                     //       .export
		.coe_f2_oe            (b22_f2_oe),                                                     //       .export
		.coe_f3_oe            (b22_f3_oe),                                                     //       .export
		.coe_f4_oe            (b22_f4_oe),                                                     //       .export
		.coe_f5_oe            (b22_f5_oe),                                                     //       .export
		.coe_f6_oe            (b22_f6_oe),                                                     //       .export
		.coe_f7_oe            (b22_f7_oe),                                                     //       .export
		.coe_f0_out           (b22_f0_out),                                                    //       .export
		.coe_f1_out           (b22_f1_out),                                                    //       .export
		.coe_f2_out           (b22_f2_out),                                                    //       .export
		.coe_f3_out           (b22_f3_out),                                                    //       .export
		.coe_f4_out           (b22_f4_out),                                                    //       .export
		.coe_f5_out           (b22_f5_out),                                                    //       .export
		.coe_f6_out           (b22_f6_out),                                                    //       .export
		.coe_f7_out           (b22_f7_out),                                                    //       .export
		.coe_f_in             (b22_f_in),                                                      //       .export
		.coe_GPIO             (b22_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b23 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b23_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b23_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b23_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b23_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b23_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b23_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b23_f1_oe),                                                     //       .export
		.coe_f2_oe            (b23_f2_oe),                                                     //       .export
		.coe_f3_oe            (b23_f3_oe),                                                     //       .export
		.coe_f4_oe            (b23_f4_oe),                                                     //       .export
		.coe_f5_oe            (b23_f5_oe),                                                     //       .export
		.coe_f6_oe            (b23_f6_oe),                                                     //       .export
		.coe_f7_oe            (b23_f7_oe),                                                     //       .export
		.coe_f0_out           (b23_f0_out),                                                    //       .export
		.coe_f1_out           (b23_f1_out),                                                    //       .export
		.coe_f2_out           (b23_f2_out),                                                    //       .export
		.coe_f3_out           (b23_f3_out),                                                    //       .export
		.coe_f4_out           (b23_f4_out),                                                    //       .export
		.coe_f5_out           (b23_f5_out),                                                    //       .export
		.coe_f6_out           (b23_f6_out),                                                    //       .export
		.coe_f7_out           (b23_f7_out),                                                    //       .export
		.coe_f_in             (b23_f_in),                                                      //       .export
		.coe_GPIO             (b23_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b24 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b24_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b24_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b24_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b24_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b24_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b24_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b24_f1_oe),                                                     //       .export
		.coe_f2_oe            (b24_f2_oe),                                                     //       .export
		.coe_f3_oe            (b24_f3_oe),                                                     //       .export
		.coe_f4_oe            (b24_f4_oe),                                                     //       .export
		.coe_f5_oe            (b24_f5_oe),                                                     //       .export
		.coe_f6_oe            (b24_f6_oe),                                                     //       .export
		.coe_f7_oe            (b24_f7_oe),                                                     //       .export
		.coe_f0_out           (b24_f0_out),                                                    //       .export
		.coe_f1_out           (b24_f1_out),                                                    //       .export
		.coe_f2_out           (b24_f2_out),                                                    //       .export
		.coe_f3_out           (b24_f3_out),                                                    //       .export
		.coe_f4_out           (b24_f4_out),                                                    //       .export
		.coe_f5_out           (b24_f5_out),                                                    //       .export
		.coe_f6_out           (b24_f6_out),                                                    //       .export
		.coe_f7_out           (b24_f7_out),                                                    //       .export
		.coe_f_in             (b24_f_in),                                                      //       .export
		.coe_GPIO             (b24_GPIO)                                                       //       .export
	);

	qsys_shield_gpioFuncSel shiled_io_b25 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                               //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                 //   MCLK.clk
		.avs_ctrl_writedata   (shiled_io_b25_ctrl_translator_avalon_anti_slave_0_writedata),   //   ctrl.writedata
		.avs_ctrl_readdata    (shiled_io_b25_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_ctrl_write       (shiled_io_b25_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_ctrl_read        (shiled_io_b25_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_ctrl_waitrequest (shiled_io_b25_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.coe_f0_oe            (b25_f0_oe),                                                     // EXPORT.export
		.coe_f1_oe            (b25_f1_oe),                                                     //       .export
		.coe_f2_oe            (b25_f2_oe),                                                     //       .export
		.coe_f3_oe            (b25_f3_oe),                                                     //       .export
		.coe_f4_oe            (b25_f4_oe),                                                     //       .export
		.coe_f5_oe            (b25_f5_oe),                                                     //       .export
		.coe_f6_oe            (b25_f6_oe),                                                     //       .export
		.coe_f7_oe            (b25_f7_oe),                                                     //       .export
		.coe_f0_out           (b25_f0_out),                                                    //       .export
		.coe_f1_out           (b25_f1_out),                                                    //       .export
		.coe_f2_out           (b25_f2_out),                                                    //       .export
		.coe_f3_out           (b25_f3_out),                                                    //       .export
		.coe_f4_out           (b25_f4_out),                                                    //       .export
		.coe_f5_out           (b25_f5_out),                                                    //       .export
		.coe_f6_out           (b25_f6_out),                                                    //       .export
		.coe_f7_out           (b25_f7_out),                                                    //       .export
		.coe_f_in             (b25_f_in),                                                      //       .export
		.coe_GPIO             (b25_GPIO)                                                       //       .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (1),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sam9_m1_translator (
		.clk                   (sam9_mclk_clk),                                              //                       clk.clk
		.reset                 (sam9_mrst_reset),                                            //                     reset.reset
		.uav_address           (sam9_m1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sam9_m1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sam9_m1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sam9_m1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sam9_m1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sam9_m1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sam9_m1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sam9_m1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sam9_m1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sam9_m1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sam9_m1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sam9_m1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sam9_m1_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (sam9_m1_byteenable),                                         //                          .byteenable
		.av_begintransfer      (sam9_m1_begintransfer),                                      //                          .begintransfer
		.av_read               (sam9_m1_read),                                               //                          .read
		.av_readdata           (sam9_m1_readdata),                                           //                          .readdata
		.av_readdatavalid      (sam9_m1_readdatavalid),                                      //                          .readdatavalid
		.av_write              (sam9_m1_write),                                              //                          .write
		.av_writedata          (sam9_m1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                       //               (terminated)
		.av_beginbursttransfer (1'b0),                                                       //               (terminated)
		.av_chipselect         (1'b0),                                                       //               (terminated)
		.av_lock               (1'b0),                                                       //               (terminated)
		.av_debugaccess        (1'b0),                                                       //               (terminated)
		.uav_clken             (),                                                           //               (terminated)
		.av_clken              (1'b1)                                                        //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_sysid_translator (
		.clk                   (sam9_mclk_clk),                                                          //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                        //                    reset.reset
		.uav_address           (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (sysid_sysid_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (sysid_sysid_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (sysid_sysid_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                       //              (terminated)
		.av_write              (),                                                                       //              (terminated)
		.av_writedata          (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_chipselect         (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) funcled_0_ledd_translator (
		.clk                   (sam9_mclk_clk),                                                             //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                           //                    reset.reset
		.uav_address           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (funcled_0_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (funcled_0_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (funcled_0_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (funcled_0_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (funcled_0_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (funcled_0_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_chipselect         (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) funcled_1_ledd_translator (
		.clk                   (sam9_mclk_clk),                                                             //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                           //                    reset.reset
		.uav_address           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (funcled_1_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (funcled_1_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (funcled_1_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (funcled_1_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (funcled_1_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (funcled_1_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_chipselect         (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) funcled_2_ledd_translator (
		.clk                   (sam9_mclk_clk),                                                             //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                           //                    reset.reset
		.uav_address           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (funcled_2_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (funcled_2_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (funcled_2_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (funcled_2_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (funcled_2_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (funcled_2_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_chipselect         (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) funcled_3_ledd_translator (
		.clk                   (sam9_mclk_clk),                                                             //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                           //                    reset.reset
		.uav_address           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (funcled_3_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (funcled_3_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (funcled_3_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (funcled_3_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (funcled_3_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (funcled_3_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_chipselect         (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shield_admin_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shield_admin_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shield_admin_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shield_admin_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shield_admin_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (shield_admin_ctrl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (shield_admin_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a0_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a0_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a0_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a0_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a0_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a0_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a1_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a1_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a1_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a1_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a1_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a1_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a2_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a2_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a2_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a2_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a2_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a2_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a3_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a3_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a3_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a3_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a3_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a3_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a4_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a4_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a4_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a4_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a4_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a4_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a5_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a5_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a5_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a5_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a5_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a5_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a6_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a6_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a6_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a6_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a6_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a6_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a7_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a7_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a7_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a7_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a7_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a7_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a8_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a8_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a8_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a8_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a8_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a8_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a9_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a9_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a9_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a9_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a9_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a9_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a10_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a10_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a10_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a10_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a10_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a10_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a11_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a11_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a11_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a11_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a11_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a11_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a13_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a13_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a13_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a13_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a13_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a13_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a12_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a12_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a12_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a12_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a12_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a12_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a14_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a14_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a14_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a14_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a14_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a14_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a15_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a15_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a15_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a15_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a15_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a15_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a17_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a17_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a17_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a17_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a17_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a17_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a16_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a16_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a16_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a16_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a16_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a16_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a18_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a18_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a18_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a18_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a18_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a18_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a19_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a19_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a19_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a19_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a19_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a19_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a20_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a20_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a20_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a20_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a20_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a20_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a21_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a21_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a21_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a21_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a21_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a21_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a22_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a22_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a22_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a22_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a22_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a22_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a23_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a23_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a23_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a23_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a23_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a23_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a24_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a24_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a24_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a24_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a24_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a24_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_a25_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_a25_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_a25_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_a25_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_a25_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_a25_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b0_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b0_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b0_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b0_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b0_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b0_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b1_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b1_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b1_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b1_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b1_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b1_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b2_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b2_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b2_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b2_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b2_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b2_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b3_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b3_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b3_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b3_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b3_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b3_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b4_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b4_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b4_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b4_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b4_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b4_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b6_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b6_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b6_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b6_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b6_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b6_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b5_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b5_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b5_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b5_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b5_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b5_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b7_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b7_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b7_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b7_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b7_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b7_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b8_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b8_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b8_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b8_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b8_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b8_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b9_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b9_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b9_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b9_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b9_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b9_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b10_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b10_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b10_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b10_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b10_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b10_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b11_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b11_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b11_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b11_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b11_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b11_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b12_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b12_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b12_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b12_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b12_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b12_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b13_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b13_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b13_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b13_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b13_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b13_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b14_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b14_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b14_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b14_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b14_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b14_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b15_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b15_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b15_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b15_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b15_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b15_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b16_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b16_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b16_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b16_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b16_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b16_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b17_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b17_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b17_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b17_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b17_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b17_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b18_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b18_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b18_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b18_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b18_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b18_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b19_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b19_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b19_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b19_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b19_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b19_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b20_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b20_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b20_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b20_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b20_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b20_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b21_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b21_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b21_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b21_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b21_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b21_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b22_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b22_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b22_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b22_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b22_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b22_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b23_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b23_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b23_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b23_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b23_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b23_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b24_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b24_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b24_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b24_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b24_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b24_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shiled_io_b25_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                 //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                               //                    reset.reset
		.uav_address           (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shiled_io_b25_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shiled_io_b25_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shiled_io_b25_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shiled_io_b25_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (shiled_io_b25_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                            //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                            //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                             //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                      //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                          //                .channel
		.rf_sink_ready           (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_004_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_004_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_004_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_004_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_004_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_004_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_005_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_005_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_005_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_005_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_005_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_005_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_006_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_006_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_006_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_006_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_006_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_006_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_007_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_007_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_007_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_007_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_007_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_007_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_008_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_008_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_008_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_008_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_008_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_008_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_009_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_009_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_009_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_009_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_009_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_009_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (92),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) funcled_0_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                       //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                     //       clk_reset.reset
		.m0_address              (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                         //                .channel
		.rf_sink_ready           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                       //       clk.clk
		.reset             (sam9_mrst_reset),                                                                     // clk_reset.reset
		.in_data           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_010_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_010_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_010_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_010_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_010_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_010_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_011_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_011_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_011_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_011_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_011_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_011_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_012_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_012_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_012_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_012_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_012_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_012_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_013_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_013_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_013_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_013_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_013_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_013_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_014_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_014_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_014_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_014_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_014_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_014_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_015_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_015_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_015_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_015_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_015_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_015_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_016_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_016_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_016_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_016_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_016_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_016_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_017_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_017_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_017_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_017_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_017_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_017_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_018_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_018_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_018_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_018_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_018_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_018_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (92),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (86),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (58),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7)
	) sam9_m1_translator_avalon_universal_master_0_agent (
		.clk              (sam9_mclk_clk),                                                       //       clk.clk
		.reset            (sam9_mrst_reset),                                                     // clk_reset.reset
		.av_address       (sam9_m1_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sam9_m1_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sam9_m1_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sam9_m1_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sam9_m1_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sam9_m1_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sam9_m1_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sam9_m1_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sam9_m1_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sam9_m1_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sam9_m1_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sam9_m1_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sam9_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sam9_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sam9_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sam9_m1_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                               //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                //          .data
		.rp_channel       (limiter_rsp_src_channel),                                             //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                       //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                         //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_019_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_019_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_019_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_019_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_019_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_019_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_020_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_020_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_020_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_020_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_020_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_020_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_021_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_021_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_021_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_021_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_021_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_021_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_022_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_022_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_022_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_022_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_022_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_022_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_023_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_023_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_023_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_023_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_023_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_023_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_024_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_024_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_024_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_024_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_024_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_024_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_025_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_025_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_025_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_025_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_025_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_025_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_026_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_026_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_026_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_026_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_026_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_026_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_027_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_027_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_027_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_027_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_027_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_027_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_028_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_028_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_028_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_028_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_028_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_028_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (92),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) funcled_1_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                       //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                     //       clk_reset.reset
		.m0_address              (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src2_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_src2_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_src2_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_src2_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src2_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src2_channel),                                                         //                .channel
		.rf_sink_ready           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                       //       clk.clk
		.reset             (sam9_mrst_reset),                                                                     // clk_reset.reset
		.in_data           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_029_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_029_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_029_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_029_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_029_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_029_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_030_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_030_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_030_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_030_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_030_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_030_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_031_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_031_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_031_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_031_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_031_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_031_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_032_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_032_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_032_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_032_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_032_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_032_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_033_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_033_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_033_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_033_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_033_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_033_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_034_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_034_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_034_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_034_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_034_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_034_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_035_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_035_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_035_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_035_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_035_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_035_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_036_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_036_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_036_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_036_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_036_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_036_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_037_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_037_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_037_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_037_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_037_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_037_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_038_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_038_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_038_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_038_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_038_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_038_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (92),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shield_admin_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src5_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_src5_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_src5_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_src5_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src5_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src5_channel),                                                            //                .channel
		.rf_sink_ready           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_039_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_039_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_039_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_039_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_039_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_039_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (92),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_sysid_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                    //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                  //       clk_reset.reset
		.m0_address              (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                      //                .channel
		.rf_sink_ready           (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                    //       clk.clk
		.reset             (sam9_mrst_reset),                                                                  // clk_reset.reset
		.in_data           (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_040_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_040_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_040_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_040_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_040_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_040_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_041_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_041_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_041_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_041_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_041_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_041_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_042_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_042_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_042_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_042_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_042_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_042_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (92),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) funcled_3_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                       //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                     //       clk_reset.reset
		.m0_address              (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src4_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_src4_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_src4_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_src4_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src4_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src4_channel),                                                         //                .channel
		.rf_sink_ready           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                       //       clk.clk
		.reset             (sam9_mrst_reset),                                                                     // clk_reset.reset
		.in_data           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_043_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_043_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_043_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_043_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_043_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_043_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_044_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_044_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_044_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_044_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_044_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_044_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_045_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_045_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_045_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_045_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_045_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_045_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_046_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_046_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_046_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_046_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_046_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_046_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_047_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_047_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_047_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_047_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_047_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_047_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_048_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_048_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_048_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_048_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_048_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_048_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (92),
		.PKT_PROTECTION_L          (92),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) funcled_2_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                       //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                     //       clk_reset.reset
		.m0_address              (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src3_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_src3_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_src3_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_src3_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src3_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src3_channel),                                                         //                .channel
		.rf_sink_ready           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                       //       clk.clk
		.reset             (sam9_mrst_reset),                                                                     // clk_reset.reset
		.in_data           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_049_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_049_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_049_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_049_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_049_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_049_source0_channel),                                                      //                .channel
		.rf_sink_ready           (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_050_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_050_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_050_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_050_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_050_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_050_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (52),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (58),
		.PKT_SRC_ID_L              (53),
		.PKT_DEST_ID_H             (64),
		.PKT_DEST_ID_L             (59),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_PROTECTION_H          (65),
		.PKT_PROTECTION_L          (65),
		.ST_CHANNEL_W              (58),
		.ST_DATA_W                 (66),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                           //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_051_source0_ready),                                                         //              cp.ready
		.cp_valid                (burst_adapter_051_source0_valid),                                                         //                .valid
		.cp_data                 (burst_adapter_051_source0_data),                                                          //                .data
		.cp_startofpacket        (burst_adapter_051_source0_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (burst_adapter_051_source0_endofpacket),                                                   //                .endofpacket
		.cp_channel              (burst_adapter_051_source0_channel),                                                       //                .channel
		.rf_sink_ready           (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (67),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                           //       clk.clk
		.reset             (sam9_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	frontier_addr_router addr_router (
		.sink_ready         (sam9_m1_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sam9_m1_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sam9_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sam9_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sam9_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                       //       clk.clk
		.reset              (sam9_mrst_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                               //       src.ready
		.src_valid          (addr_router_src_valid),                                               //          .valid
		.src_data           (addr_router_src_data),                                                //          .data
		.src_channel        (addr_router_src_channel),                                             //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                          //          .endofpacket
	);

	frontier_id_router id_router (
		.sink_ready         (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                          //       clk.clk
		.reset              (sam9_mrst_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                    //       src.ready
		.src_valid          (id_router_src_valid),                                                    //          .valid
		.src_data           (id_router_src_data),                                                     //          .data
		.src_channel        (id_router_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                               //          .endofpacket
	);

	frontier_id_router id_router_001 (
		.sink_ready         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                             //       clk.clk
		.reset              (sam9_mrst_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                   //       src.ready
		.src_valid          (id_router_001_src_valid),                                                   //          .valid
		.src_data           (id_router_001_src_data),                                                    //          .data
		.src_channel        (id_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                              //          .endofpacket
	);

	frontier_id_router id_router_002 (
		.sink_ready         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                             //       clk.clk
		.reset              (sam9_mrst_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                   //       src.ready
		.src_valid          (id_router_002_src_valid),                                                   //          .valid
		.src_data           (id_router_002_src_data),                                                    //          .data
		.src_channel        (id_router_002_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                              //          .endofpacket
	);

	frontier_id_router id_router_003 (
		.sink_ready         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                             //       clk.clk
		.reset              (sam9_mrst_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                   //       src.ready
		.src_valid          (id_router_003_src_valid),                                                   //          .valid
		.src_data           (id_router_003_src_data),                                                    //          .data
		.src_channel        (id_router_003_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                              //          .endofpacket
	);

	frontier_id_router id_router_004 (
		.sink_ready         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                             //       clk.clk
		.reset              (sam9_mrst_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                   //       src.ready
		.src_valid          (id_router_004_src_valid),                                                   //          .valid
		.src_data           (id_router_004_src_data),                                                    //          .data
		.src_channel        (id_router_004_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                              //          .endofpacket
	);

	frontier_id_router id_router_005 (
		.sink_ready         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                      //       src.ready
		.src_valid          (id_router_005_src_valid),                                                      //          .valid
		.src_data           (id_router_005_src_data),                                                       //          .data
		.src_channel        (id_router_005_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_006 (
		.sink_ready         (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                      //       src.ready
		.src_valid          (id_router_006_src_valid),                                                      //          .valid
		.src_data           (id_router_006_src_data),                                                       //          .data
		.src_channel        (id_router_006_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_007 (
		.sink_ready         (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a1_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                      //       src.ready
		.src_valid          (id_router_007_src_valid),                                                      //          .valid
		.src_data           (id_router_007_src_data),                                                       //          .data
		.src_channel        (id_router_007_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_008 (
		.sink_ready         (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a2_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                      //       src.ready
		.src_valid          (id_router_008_src_valid),                                                      //          .valid
		.src_data           (id_router_008_src_data),                                                       //          .data
		.src_channel        (id_router_008_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_009 (
		.sink_ready         (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a3_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                      //       src.ready
		.src_valid          (id_router_009_src_valid),                                                      //          .valid
		.src_data           (id_router_009_src_data),                                                       //          .data
		.src_channel        (id_router_009_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_010 (
		.sink_ready         (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a4_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                      //       src.ready
		.src_valid          (id_router_010_src_valid),                                                      //          .valid
		.src_data           (id_router_010_src_data),                                                       //          .data
		.src_channel        (id_router_010_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_011 (
		.sink_ready         (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a5_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                      //       src.ready
		.src_valid          (id_router_011_src_valid),                                                      //          .valid
		.src_data           (id_router_011_src_data),                                                       //          .data
		.src_channel        (id_router_011_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_012 (
		.sink_ready         (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a6_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                      //       src.ready
		.src_valid          (id_router_012_src_valid),                                                      //          .valid
		.src_data           (id_router_012_src_data),                                                       //          .data
		.src_channel        (id_router_012_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_013 (
		.sink_ready         (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a7_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                      //       src.ready
		.src_valid          (id_router_013_src_valid),                                                      //          .valid
		.src_data           (id_router_013_src_data),                                                       //          .data
		.src_channel        (id_router_013_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_014 (
		.sink_ready         (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a8_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                      //       src.ready
		.src_valid          (id_router_014_src_valid),                                                      //          .valid
		.src_data           (id_router_014_src_data),                                                       //          .data
		.src_channel        (id_router_014_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_015 (
		.sink_ready         (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a9_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                      //       src.ready
		.src_valid          (id_router_015_src_valid),                                                      //          .valid
		.src_data           (id_router_015_src_data),                                                       //          .data
		.src_channel        (id_router_015_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_016 (
		.sink_ready         (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a10_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                       //       src.ready
		.src_valid          (id_router_016_src_valid),                                                       //          .valid
		.src_data           (id_router_016_src_data),                                                        //          .data
		.src_channel        (id_router_016_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_017 (
		.sink_ready         (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a11_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                       //       src.ready
		.src_valid          (id_router_017_src_valid),                                                       //          .valid
		.src_data           (id_router_017_src_data),                                                        //          .data
		.src_channel        (id_router_017_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_018 (
		.sink_ready         (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a13_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                       //       src.ready
		.src_valid          (id_router_018_src_valid),                                                       //          .valid
		.src_data           (id_router_018_src_data),                                                        //          .data
		.src_channel        (id_router_018_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_019 (
		.sink_ready         (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a12_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                       //       src.ready
		.src_valid          (id_router_019_src_valid),                                                       //          .valid
		.src_data           (id_router_019_src_data),                                                        //          .data
		.src_channel        (id_router_019_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_020 (
		.sink_ready         (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a14_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                       //       src.ready
		.src_valid          (id_router_020_src_valid),                                                       //          .valid
		.src_data           (id_router_020_src_data),                                                        //          .data
		.src_channel        (id_router_020_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_021 (
		.sink_ready         (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a15_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                                       //       src.ready
		.src_valid          (id_router_021_src_valid),                                                       //          .valid
		.src_data           (id_router_021_src_data),                                                        //          .data
		.src_channel        (id_router_021_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_022 (
		.sink_ready         (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a17_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                                       //       src.ready
		.src_valid          (id_router_022_src_valid),                                                       //          .valid
		.src_data           (id_router_022_src_data),                                                        //          .data
		.src_channel        (id_router_022_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_023 (
		.sink_ready         (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a16_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                                       //       src.ready
		.src_valid          (id_router_023_src_valid),                                                       //          .valid
		.src_data           (id_router_023_src_data),                                                        //          .data
		.src_channel        (id_router_023_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_024 (
		.sink_ready         (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a18_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                                       //       src.ready
		.src_valid          (id_router_024_src_valid),                                                       //          .valid
		.src_data           (id_router_024_src_data),                                                        //          .data
		.src_channel        (id_router_024_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_025 (
		.sink_ready         (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a19_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                                       //       src.ready
		.src_valid          (id_router_025_src_valid),                                                       //          .valid
		.src_data           (id_router_025_src_data),                                                        //          .data
		.src_channel        (id_router_025_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_026 (
		.sink_ready         (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a20_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_026_src_ready),                                                       //       src.ready
		.src_valid          (id_router_026_src_valid),                                                       //          .valid
		.src_data           (id_router_026_src_data),                                                        //          .data
		.src_channel        (id_router_026_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_026_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_026_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_027 (
		.sink_ready         (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a21_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_027_src_ready),                                                       //       src.ready
		.src_valid          (id_router_027_src_valid),                                                       //          .valid
		.src_data           (id_router_027_src_data),                                                        //          .data
		.src_channel        (id_router_027_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_027_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_027_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_028 (
		.sink_ready         (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a22_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_028_src_ready),                                                       //       src.ready
		.src_valid          (id_router_028_src_valid),                                                       //          .valid
		.src_data           (id_router_028_src_data),                                                        //          .data
		.src_channel        (id_router_028_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_028_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_028_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_029 (
		.sink_ready         (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a23_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_029_src_ready),                                                       //       src.ready
		.src_valid          (id_router_029_src_valid),                                                       //          .valid
		.src_data           (id_router_029_src_data),                                                        //          .data
		.src_channel        (id_router_029_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_029_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_029_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_030 (
		.sink_ready         (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a24_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_030_src_ready),                                                       //       src.ready
		.src_valid          (id_router_030_src_valid),                                                       //          .valid
		.src_data           (id_router_030_src_data),                                                        //          .data
		.src_channel        (id_router_030_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_030_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_030_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_031 (
		.sink_ready         (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_a25_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_031_src_ready),                                                       //       src.ready
		.src_valid          (id_router_031_src_valid),                                                       //          .valid
		.src_data           (id_router_031_src_data),                                                        //          .data
		.src_channel        (id_router_031_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_031_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_031_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_032 (
		.sink_ready         (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_032_src_ready),                                                      //       src.ready
		.src_valid          (id_router_032_src_valid),                                                      //          .valid
		.src_data           (id_router_032_src_data),                                                       //          .data
		.src_channel        (id_router_032_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_032_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_032_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_033 (
		.sink_ready         (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b1_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_033_src_ready),                                                      //       src.ready
		.src_valid          (id_router_033_src_valid),                                                      //          .valid
		.src_data           (id_router_033_src_data),                                                       //          .data
		.src_channel        (id_router_033_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_033_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_033_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_034 (
		.sink_ready         (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b2_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_034_src_ready),                                                      //       src.ready
		.src_valid          (id_router_034_src_valid),                                                      //          .valid
		.src_data           (id_router_034_src_data),                                                       //          .data
		.src_channel        (id_router_034_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_034_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_034_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_035 (
		.sink_ready         (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b3_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_035_src_ready),                                                      //       src.ready
		.src_valid          (id_router_035_src_valid),                                                      //          .valid
		.src_data           (id_router_035_src_data),                                                       //          .data
		.src_channel        (id_router_035_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_035_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_035_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_036 (
		.sink_ready         (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b4_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_036_src_ready),                                                      //       src.ready
		.src_valid          (id_router_036_src_valid),                                                      //          .valid
		.src_data           (id_router_036_src_data),                                                       //          .data
		.src_channel        (id_router_036_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_036_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_036_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_037 (
		.sink_ready         (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b6_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_037_src_ready),                                                      //       src.ready
		.src_valid          (id_router_037_src_valid),                                                      //          .valid
		.src_data           (id_router_037_src_data),                                                       //          .data
		.src_channel        (id_router_037_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_037_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_037_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_038 (
		.sink_ready         (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b5_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_038_src_ready),                                                      //       src.ready
		.src_valid          (id_router_038_src_valid),                                                      //          .valid
		.src_data           (id_router_038_src_data),                                                       //          .data
		.src_channel        (id_router_038_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_038_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_038_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_039 (
		.sink_ready         (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b7_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_039_src_ready),                                                      //       src.ready
		.src_valid          (id_router_039_src_valid),                                                      //          .valid
		.src_data           (id_router_039_src_data),                                                       //          .data
		.src_channel        (id_router_039_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_039_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_039_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_040 (
		.sink_ready         (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b8_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_040_src_ready),                                                      //       src.ready
		.src_valid          (id_router_040_src_valid),                                                      //          .valid
		.src_data           (id_router_040_src_data),                                                       //          .data
		.src_channel        (id_router_040_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_040_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_040_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_041 (
		.sink_ready         (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b9_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_041_src_ready),                                                      //       src.ready
		.src_valid          (id_router_041_src_valid),                                                      //          .valid
		.src_data           (id_router_041_src_data),                                                       //          .data
		.src_channel        (id_router_041_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_041_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_041_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router_006 id_router_042 (
		.sink_ready         (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b10_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_042_src_ready),                                                       //       src.ready
		.src_valid          (id_router_042_src_valid),                                                       //          .valid
		.src_data           (id_router_042_src_data),                                                        //          .data
		.src_channel        (id_router_042_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_042_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_042_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_043 (
		.sink_ready         (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b11_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_043_src_ready),                                                       //       src.ready
		.src_valid          (id_router_043_src_valid),                                                       //          .valid
		.src_data           (id_router_043_src_data),                                                        //          .data
		.src_channel        (id_router_043_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_043_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_043_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_044 (
		.sink_ready         (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b12_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_044_src_ready),                                                       //       src.ready
		.src_valid          (id_router_044_src_valid),                                                       //          .valid
		.src_data           (id_router_044_src_data),                                                        //          .data
		.src_channel        (id_router_044_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_044_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_044_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_045 (
		.sink_ready         (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b13_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_045_src_ready),                                                       //       src.ready
		.src_valid          (id_router_045_src_valid),                                                       //          .valid
		.src_data           (id_router_045_src_data),                                                        //          .data
		.src_channel        (id_router_045_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_045_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_045_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_046 (
		.sink_ready         (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b14_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_046_src_ready),                                                       //       src.ready
		.src_valid          (id_router_046_src_valid),                                                       //          .valid
		.src_data           (id_router_046_src_data),                                                        //          .data
		.src_channel        (id_router_046_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_046_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_046_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_047 (
		.sink_ready         (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b15_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_047_src_ready),                                                       //       src.ready
		.src_valid          (id_router_047_src_valid),                                                       //          .valid
		.src_data           (id_router_047_src_data),                                                        //          .data
		.src_channel        (id_router_047_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_047_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_047_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_048 (
		.sink_ready         (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b16_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_048_src_ready),                                                       //       src.ready
		.src_valid          (id_router_048_src_valid),                                                       //          .valid
		.src_data           (id_router_048_src_data),                                                        //          .data
		.src_channel        (id_router_048_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_048_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_048_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_049 (
		.sink_ready         (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b17_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_049_src_ready),                                                       //       src.ready
		.src_valid          (id_router_049_src_valid),                                                       //          .valid
		.src_data           (id_router_049_src_data),                                                        //          .data
		.src_channel        (id_router_049_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_049_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_049_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_050 (
		.sink_ready         (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b18_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_050_src_ready),                                                       //       src.ready
		.src_valid          (id_router_050_src_valid),                                                       //          .valid
		.src_data           (id_router_050_src_data),                                                        //          .data
		.src_channel        (id_router_050_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_050_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_050_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_051 (
		.sink_ready         (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b19_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_051_src_ready),                                                       //       src.ready
		.src_valid          (id_router_051_src_valid),                                                       //          .valid
		.src_data           (id_router_051_src_data),                                                        //          .data
		.src_channel        (id_router_051_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_051_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_051_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_052 (
		.sink_ready         (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b20_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_052_src_ready),                                                       //       src.ready
		.src_valid          (id_router_052_src_valid),                                                       //          .valid
		.src_data           (id_router_052_src_data),                                                        //          .data
		.src_channel        (id_router_052_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_052_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_052_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_053 (
		.sink_ready         (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b21_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_053_src_ready),                                                       //       src.ready
		.src_valid          (id_router_053_src_valid),                                                       //          .valid
		.src_data           (id_router_053_src_data),                                                        //          .data
		.src_channel        (id_router_053_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_053_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_053_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_054 (
		.sink_ready         (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b22_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_054_src_ready),                                                       //       src.ready
		.src_valid          (id_router_054_src_valid),                                                       //          .valid
		.src_data           (id_router_054_src_data),                                                        //          .data
		.src_channel        (id_router_054_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_054_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_054_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_055 (
		.sink_ready         (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b23_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_055_src_ready),                                                       //       src.ready
		.src_valid          (id_router_055_src_valid),                                                       //          .valid
		.src_data           (id_router_055_src_data),                                                        //          .data
		.src_channel        (id_router_055_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_055_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_055_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_056 (
		.sink_ready         (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b24_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_056_src_ready),                                                       //       src.ready
		.src_valid          (id_router_056_src_valid),                                                       //          .valid
		.src_data           (id_router_056_src_data),                                                        //          .data
		.src_channel        (id_router_056_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_056_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_056_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router_006 id_router_057 (
		.sink_ready         (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shiled_io_b25_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                 //       clk.clk
		.reset              (sam9_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_057_src_ready),                                                       //       src.ready
		.src_valid          (id_router_057_src_valid),                                                       //          .valid
		.src_data           (id_router_057_src_data),                                                        //          .data
		.src_channel        (id_router_057_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_057_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_057_src_endofpacket)                                                  //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (86),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (3),
		.PIPELINED                 (0),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (58),
		.VALID_WIDTH               (58),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (sam9_mclk_clk),                  //       clk.clk
		.reset                  (sam9_mrst_reset),                // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter (
		.clk                   (sam9_mclk_clk),                       //       cr0.clk
		.reset                 (sam9_mrst_reset),                     // cr0_reset.reset
		.sink0_valid           (width_adapter_052_src_valid),         //     sink0.valid
		.sink0_data            (width_adapter_052_src_data),          //          .data
		.sink0_channel         (width_adapter_052_src_channel),       //          .channel
		.sink0_startofpacket   (width_adapter_052_src_startofpacket), //          .startofpacket
		.sink0_endofpacket     (width_adapter_052_src_endofpacket),   //          .endofpacket
		.sink0_ready           (width_adapter_052_src_ready),         //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_001 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_056_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_056_src_data),              //          .data
		.sink0_channel         (width_adapter_056_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_056_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_056_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_056_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_002 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_026_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_026_src_data),              //          .data
		.sink0_channel         (width_adapter_026_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_026_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_026_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_026_src_ready),             //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_003 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_022_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_022_src_data),              //          .data
		.sink0_channel         (width_adapter_022_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_022_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_022_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_022_src_ready),             //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_004 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_004_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_004_source0_data),          //          .data
		.source0_channel       (burst_adapter_004_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_004_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_004_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_004_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_005 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),                 //     sink0.valid
		.sink0_data            (width_adapter_src_data),                  //          .data
		.sink0_channel         (width_adapter_src_channel),               //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),         //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),           //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),                 //          .ready
		.source0_valid         (burst_adapter_005_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_005_source0_data),          //          .data
		.source0_channel       (burst_adapter_005_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_005_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_005_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_005_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_006 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_090_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_090_src_data),              //          .data
		.sink0_channel         (width_adapter_090_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_090_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_090_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_090_src_ready),             //          .ready
		.source0_valid         (burst_adapter_006_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_006_source0_data),          //          .data
		.source0_channel       (burst_adapter_006_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_006_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_006_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_006_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_007 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_020_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_020_src_data),              //          .data
		.sink0_channel         (width_adapter_020_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_020_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_020_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_020_src_ready),             //          .ready
		.source0_valid         (burst_adapter_007_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_007_source0_data),          //          .data
		.source0_channel       (burst_adapter_007_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_007_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_007_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_007_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_008 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_038_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_038_src_data),              //          .data
		.sink0_channel         (width_adapter_038_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_038_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_038_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_038_src_ready),             //          .ready
		.source0_valid         (burst_adapter_008_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_008_source0_data),          //          .data
		.source0_channel       (burst_adapter_008_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_008_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_008_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_008_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_009 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_054_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_054_src_data),              //          .data
		.sink0_channel         (width_adapter_054_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_054_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_054_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_054_src_ready),             //          .ready
		.source0_valid         (burst_adapter_009_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_009_source0_data),          //          .data
		.source0_channel       (burst_adapter_009_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_009_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_009_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_009_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_010 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_012_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_012_src_data),              //          .data
		.sink0_channel         (width_adapter_012_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_012_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_012_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_012_src_ready),             //          .ready
		.source0_valid         (burst_adapter_010_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_010_source0_data),          //          .data
		.source0_channel       (burst_adapter_010_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_010_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_010_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_010_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_011 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_008_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_008_src_data),              //          .data
		.sink0_channel         (width_adapter_008_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_008_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_008_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_008_src_ready),             //          .ready
		.source0_valid         (burst_adapter_011_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_011_source0_data),          //          .data
		.source0_channel       (burst_adapter_011_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_011_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_011_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_011_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_012 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_040_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_040_src_data),              //          .data
		.sink0_channel         (width_adapter_040_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_040_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_040_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_040_src_ready),             //          .ready
		.source0_valid         (burst_adapter_012_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_012_source0_data),          //          .data
		.source0_channel       (burst_adapter_012_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_012_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_012_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_012_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_013 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_074_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_074_src_data),              //          .data
		.sink0_channel         (width_adapter_074_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_074_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_074_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_074_src_ready),             //          .ready
		.source0_valid         (burst_adapter_013_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_013_source0_data),          //          .data
		.source0_channel       (burst_adapter_013_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_013_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_013_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_013_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_014 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_032_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_032_src_data),              //          .data
		.sink0_channel         (width_adapter_032_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_032_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_032_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_032_src_ready),             //          .ready
		.source0_valid         (burst_adapter_014_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_014_source0_data),          //          .data
		.source0_channel       (burst_adapter_014_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_014_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_014_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_014_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_015 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_068_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_068_src_data),              //          .data
		.sink0_channel         (width_adapter_068_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_068_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_068_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_068_src_ready),             //          .ready
		.source0_valid         (burst_adapter_015_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_015_source0_data),          //          .data
		.source0_channel       (burst_adapter_015_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_015_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_015_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_015_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_016 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_100_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_100_src_data),              //          .data
		.sink0_channel         (width_adapter_100_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_100_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_100_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_100_src_ready),             //          .ready
		.source0_valid         (burst_adapter_016_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_016_source0_data),          //          .data
		.source0_channel       (burst_adapter_016_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_016_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_016_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_016_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_017 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_066_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_066_src_data),              //          .data
		.sink0_channel         (width_adapter_066_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_066_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_066_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_066_src_ready),             //          .ready
		.source0_valid         (burst_adapter_017_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_017_source0_data),          //          .data
		.source0_channel       (burst_adapter_017_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_017_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_017_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_017_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_018 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_092_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_092_src_data),              //          .data
		.sink0_channel         (width_adapter_092_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_092_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_092_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_092_src_ready),             //          .ready
		.source0_valid         (burst_adapter_018_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_018_source0_data),          //          .data
		.source0_channel       (burst_adapter_018_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_018_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_018_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_018_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_019 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_048_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_048_src_data),              //          .data
		.sink0_channel         (width_adapter_048_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_048_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_048_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_048_src_ready),             //          .ready
		.source0_valid         (burst_adapter_019_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_019_source0_data),          //          .data
		.source0_channel       (burst_adapter_019_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_019_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_019_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_019_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_020 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_084_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_084_src_data),              //          .data
		.sink0_channel         (width_adapter_084_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_084_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_084_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_084_src_ready),             //          .ready
		.source0_valid         (burst_adapter_020_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_020_source0_data),          //          .data
		.source0_channel       (burst_adapter_020_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_020_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_020_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_020_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_021 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_050_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_050_src_data),              //          .data
		.sink0_channel         (width_adapter_050_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_050_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_050_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_050_src_ready),             //          .ready
		.source0_valid         (burst_adapter_021_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_021_source0_data),          //          .data
		.source0_channel       (burst_adapter_021_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_021_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_021_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_021_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_022 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_082_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_082_src_data),              //          .data
		.sink0_channel         (width_adapter_082_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_082_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_082_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_082_src_ready),             //          .ready
		.source0_valid         (burst_adapter_022_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_022_source0_data),          //          .data
		.source0_channel       (burst_adapter_022_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_022_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_022_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_022_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_023 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_014_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_014_src_data),              //          .data
		.sink0_channel         (width_adapter_014_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_014_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_014_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_014_src_ready),             //          .ready
		.source0_valid         (burst_adapter_023_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_023_source0_data),          //          .data
		.source0_channel       (burst_adapter_023_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_023_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_023_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_023_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_024 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_094_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_094_src_data),              //          .data
		.sink0_channel         (width_adapter_094_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_094_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_094_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_094_src_ready),             //          .ready
		.source0_valid         (burst_adapter_024_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_024_source0_data),          //          .data
		.source0_channel       (burst_adapter_024_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_024_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_024_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_024_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_025 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_006_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_006_src_data),              //          .data
		.sink0_channel         (width_adapter_006_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_006_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_006_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_006_src_ready),             //          .ready
		.source0_valid         (burst_adapter_025_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_025_source0_data),          //          .data
		.source0_channel       (burst_adapter_025_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_025_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_025_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_025_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_026 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_064_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_064_src_data),              //          .data
		.sink0_channel         (width_adapter_064_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_064_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_064_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_064_src_ready),             //          .ready
		.source0_valid         (burst_adapter_026_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_026_source0_data),          //          .data
		.source0_channel       (burst_adapter_026_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_026_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_026_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_026_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_027 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_028_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_028_src_data),              //          .data
		.sink0_channel         (width_adapter_028_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_028_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_028_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_028_src_ready),             //          .ready
		.source0_valid         (burst_adapter_027_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_027_source0_data),          //          .data
		.source0_channel       (burst_adapter_027_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_027_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_027_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_027_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_028 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_072_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_072_src_data),              //          .data
		.sink0_channel         (width_adapter_072_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_072_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_072_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_072_src_ready),             //          .ready
		.source0_valid         (burst_adapter_028_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_028_source0_data),          //          .data
		.source0_channel       (burst_adapter_028_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_028_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_028_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_028_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_029 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_076_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_076_src_data),              //          .data
		.sink0_channel         (width_adapter_076_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_076_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_076_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_076_src_ready),             //          .ready
		.source0_valid         (burst_adapter_029_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_029_source0_data),          //          .data
		.source0_channel       (burst_adapter_029_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_029_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_029_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_029_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_030 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_080_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_080_src_data),              //          .data
		.sink0_channel         (width_adapter_080_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_080_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_080_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_080_src_ready),             //          .ready
		.source0_valid         (burst_adapter_030_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_030_source0_data),          //          .data
		.source0_channel       (burst_adapter_030_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_030_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_030_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_030_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_031 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_062_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_062_src_data),              //          .data
		.sink0_channel         (width_adapter_062_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_062_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_062_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_062_src_ready),             //          .ready
		.source0_valid         (burst_adapter_031_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_031_source0_data),          //          .data
		.source0_channel       (burst_adapter_031_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_031_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_031_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_031_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_032 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_070_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_070_src_data),              //          .data
		.sink0_channel         (width_adapter_070_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_070_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_070_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_070_src_ready),             //          .ready
		.source0_valid         (burst_adapter_032_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_032_source0_data),          //          .data
		.source0_channel       (burst_adapter_032_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_032_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_032_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_032_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_033 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_044_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_044_src_data),              //          .data
		.sink0_channel         (width_adapter_044_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_044_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_044_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_044_src_ready),             //          .ready
		.source0_valid         (burst_adapter_033_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_033_source0_data),          //          .data
		.source0_channel       (burst_adapter_033_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_033_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_033_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_033_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_034 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_098_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_098_src_data),              //          .data
		.sink0_channel         (width_adapter_098_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_098_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_098_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_098_src_ready),             //          .ready
		.source0_valid         (burst_adapter_034_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_034_source0_data),          //          .data
		.source0_channel       (burst_adapter_034_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_034_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_034_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_034_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_035 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_078_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_078_src_data),              //          .data
		.sink0_channel         (width_adapter_078_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_078_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_078_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_078_src_ready),             //          .ready
		.source0_valid         (burst_adapter_035_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_035_source0_data),          //          .data
		.source0_channel       (burst_adapter_035_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_035_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_035_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_035_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_036 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_102_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_102_src_data),              //          .data
		.sink0_channel         (width_adapter_102_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_102_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_102_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_102_src_ready),             //          .ready
		.source0_valid         (burst_adapter_036_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_036_source0_data),          //          .data
		.source0_channel       (burst_adapter_036_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_036_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_036_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_036_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_037 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_042_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_042_src_data),              //          .data
		.sink0_channel         (width_adapter_042_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_042_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_042_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_042_src_ready),             //          .ready
		.source0_valid         (burst_adapter_037_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_037_source0_data),          //          .data
		.source0_channel       (burst_adapter_037_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_037_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_037_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_037_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_038 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_088_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_088_src_data),              //          .data
		.sink0_channel         (width_adapter_088_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_088_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_088_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_088_src_ready),             //          .ready
		.source0_valid         (burst_adapter_038_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_038_source0_data),          //          .data
		.source0_channel       (burst_adapter_038_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_038_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_038_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_038_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_039 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_096_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_096_src_data),              //          .data
		.sink0_channel         (width_adapter_096_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_096_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_096_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_096_src_ready),             //          .ready
		.source0_valid         (burst_adapter_039_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_039_source0_data),          //          .data
		.source0_channel       (burst_adapter_039_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_039_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_039_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_039_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_040 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_030_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_030_src_data),              //          .data
		.sink0_channel         (width_adapter_030_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_030_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_030_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_030_src_ready),             //          .ready
		.source0_valid         (burst_adapter_040_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_040_source0_data),          //          .data
		.source0_channel       (burst_adapter_040_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_040_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_040_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_040_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_041 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_060_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_060_src_data),              //          .data
		.sink0_channel         (width_adapter_060_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_060_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_060_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_060_src_ready),             //          .ready
		.source0_valid         (burst_adapter_041_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_041_source0_data),          //          .data
		.source0_channel       (burst_adapter_041_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_041_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_041_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_041_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_042 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_018_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_018_src_data),              //          .data
		.sink0_channel         (width_adapter_018_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_018_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_018_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_018_src_ready),             //          .ready
		.source0_valid         (burst_adapter_042_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_042_source0_data),          //          .data
		.source0_channel       (burst_adapter_042_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_042_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_042_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_042_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_043 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_016_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_016_src_data),              //          .data
		.sink0_channel         (width_adapter_016_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_016_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_016_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_016_src_ready),             //          .ready
		.source0_valid         (burst_adapter_043_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_043_source0_data),          //          .data
		.source0_channel       (burst_adapter_043_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_043_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_043_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_043_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_044 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_058_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_058_src_data),              //          .data
		.sink0_channel         (width_adapter_058_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_058_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_058_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_058_src_ready),             //          .ready
		.source0_valid         (burst_adapter_044_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_044_source0_data),          //          .data
		.source0_channel       (burst_adapter_044_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_044_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_044_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_044_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_045 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_086_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_086_src_data),              //          .data
		.sink0_channel         (width_adapter_086_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_086_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_086_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_086_src_ready),             //          .ready
		.source0_valid         (burst_adapter_045_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_045_source0_data),          //          .data
		.source0_channel       (burst_adapter_045_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_045_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_045_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_045_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_046 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_024_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_024_src_data),              //          .data
		.sink0_channel         (width_adapter_024_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_024_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_024_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_024_src_ready),             //          .ready
		.source0_valid         (burst_adapter_046_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_046_source0_data),          //          .data
		.source0_channel       (burst_adapter_046_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_046_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_046_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_046_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_047 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_034_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_034_src_data),              //          .data
		.sink0_channel         (width_adapter_034_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_034_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_034_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_034_src_ready),             //          .ready
		.source0_valid         (burst_adapter_047_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_047_source0_data),          //          .data
		.source0_channel       (burst_adapter_047_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_047_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_047_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_047_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_048 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_048_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_048_source0_data),          //          .data
		.source0_channel       (burst_adapter_048_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_048_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_048_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_048_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_049 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_010_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_010_src_data),              //          .data
		.sink0_channel         (width_adapter_010_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_010_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_010_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_010_src_ready),             //          .ready
		.source0_valid         (burst_adapter_049_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_049_source0_data),          //          .data
		.source0_channel       (burst_adapter_049_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_049_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_049_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_049_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_050 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_046_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_046_src_data),              //          .data
		.sink0_channel         (width_adapter_046_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_046_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_046_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_046_src_ready),             //          .ready
		.source0_valid         (burst_adapter_050_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_050_source0_data),          //          .data
		.source0_channel       (burst_adapter_050_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_050_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_050_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_050_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (52),
		.PKT_BYTE_CNT_H            (48),
		.PKT_BYTE_CNT_L            (46),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURSTWRAP_H           (51),
		.PKT_BURSTWRAP_L           (49),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.ST_DATA_W                 (66),
		.ST_CHANNEL_W              (58),
		.OUT_BYTE_CNT_H            (46),
		.OUT_BURSTWRAP_H           (51),
		.COMPRESSED_READ_SUPPORT   (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_051 (
		.clk                   (sam9_mclk_clk),                           //       cr0.clk
		.reset                 (sam9_mrst_reset),                         // cr0_reset.reset
		.sink0_valid           (width_adapter_036_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_036_src_data),              //          .data
		.sink0_channel         (width_adapter_036_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_036_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_036_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_036_src_ready),             //          .ready
		.source0_valid         (burst_adapter_051_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_051_source0_data),          //          .data
		.source0_channel       (burst_adapter_051_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_051_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_051_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_051_source0_ready)          //          .ready
	);

	frontier_cmd_xbar_demux cmd_xbar_demux (
		.clk                 (sam9_mclk_clk),                      //        clk.clk
		.reset               (sam9_mrst_reset),                    //  clk_reset.reset
		.sink_ready          (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_cmd_src_channel),            //           .channel
		.sink_data           (limiter_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_src17_endofpacket),   //           .endofpacket
		.src18_ready         (cmd_xbar_demux_src18_ready),         //      src18.ready
		.src18_valid         (cmd_xbar_demux_src18_valid),         //           .valid
		.src18_data          (cmd_xbar_demux_src18_data),          //           .data
		.src18_channel       (cmd_xbar_demux_src18_channel),       //           .channel
		.src18_startofpacket (cmd_xbar_demux_src18_startofpacket), //           .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_src18_endofpacket),   //           .endofpacket
		.src19_ready         (cmd_xbar_demux_src19_ready),         //      src19.ready
		.src19_valid         (cmd_xbar_demux_src19_valid),         //           .valid
		.src19_data          (cmd_xbar_demux_src19_data),          //           .data
		.src19_channel       (cmd_xbar_demux_src19_channel),       //           .channel
		.src19_startofpacket (cmd_xbar_demux_src19_startofpacket), //           .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_src19_endofpacket),   //           .endofpacket
		.src20_ready         (cmd_xbar_demux_src20_ready),         //      src20.ready
		.src20_valid         (cmd_xbar_demux_src20_valid),         //           .valid
		.src20_data          (cmd_xbar_demux_src20_data),          //           .data
		.src20_channel       (cmd_xbar_demux_src20_channel),       //           .channel
		.src20_startofpacket (cmd_xbar_demux_src20_startofpacket), //           .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_src20_endofpacket),   //           .endofpacket
		.src21_ready         (cmd_xbar_demux_src21_ready),         //      src21.ready
		.src21_valid         (cmd_xbar_demux_src21_valid),         //           .valid
		.src21_data          (cmd_xbar_demux_src21_data),          //           .data
		.src21_channel       (cmd_xbar_demux_src21_channel),       //           .channel
		.src21_startofpacket (cmd_xbar_demux_src21_startofpacket), //           .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_src21_endofpacket),   //           .endofpacket
		.src22_ready         (cmd_xbar_demux_src22_ready),         //      src22.ready
		.src22_valid         (cmd_xbar_demux_src22_valid),         //           .valid
		.src22_data          (cmd_xbar_demux_src22_data),          //           .data
		.src22_channel       (cmd_xbar_demux_src22_channel),       //           .channel
		.src22_startofpacket (cmd_xbar_demux_src22_startofpacket), //           .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_src22_endofpacket),   //           .endofpacket
		.src23_ready         (cmd_xbar_demux_src23_ready),         //      src23.ready
		.src23_valid         (cmd_xbar_demux_src23_valid),         //           .valid
		.src23_data          (cmd_xbar_demux_src23_data),          //           .data
		.src23_channel       (cmd_xbar_demux_src23_channel),       //           .channel
		.src23_startofpacket (cmd_xbar_demux_src23_startofpacket), //           .startofpacket
		.src23_endofpacket   (cmd_xbar_demux_src23_endofpacket),   //           .endofpacket
		.src24_ready         (cmd_xbar_demux_src24_ready),         //      src24.ready
		.src24_valid         (cmd_xbar_demux_src24_valid),         //           .valid
		.src24_data          (cmd_xbar_demux_src24_data),          //           .data
		.src24_channel       (cmd_xbar_demux_src24_channel),       //           .channel
		.src24_startofpacket (cmd_xbar_demux_src24_startofpacket), //           .startofpacket
		.src24_endofpacket   (cmd_xbar_demux_src24_endofpacket),   //           .endofpacket
		.src25_ready         (cmd_xbar_demux_src25_ready),         //      src25.ready
		.src25_valid         (cmd_xbar_demux_src25_valid),         //           .valid
		.src25_data          (cmd_xbar_demux_src25_data),          //           .data
		.src25_channel       (cmd_xbar_demux_src25_channel),       //           .channel
		.src25_startofpacket (cmd_xbar_demux_src25_startofpacket), //           .startofpacket
		.src25_endofpacket   (cmd_xbar_demux_src25_endofpacket),   //           .endofpacket
		.src26_ready         (cmd_xbar_demux_src26_ready),         //      src26.ready
		.src26_valid         (cmd_xbar_demux_src26_valid),         //           .valid
		.src26_data          (cmd_xbar_demux_src26_data),          //           .data
		.src26_channel       (cmd_xbar_demux_src26_channel),       //           .channel
		.src26_startofpacket (cmd_xbar_demux_src26_startofpacket), //           .startofpacket
		.src26_endofpacket   (cmd_xbar_demux_src26_endofpacket),   //           .endofpacket
		.src27_ready         (cmd_xbar_demux_src27_ready),         //      src27.ready
		.src27_valid         (cmd_xbar_demux_src27_valid),         //           .valid
		.src27_data          (cmd_xbar_demux_src27_data),          //           .data
		.src27_channel       (cmd_xbar_demux_src27_channel),       //           .channel
		.src27_startofpacket (cmd_xbar_demux_src27_startofpacket), //           .startofpacket
		.src27_endofpacket   (cmd_xbar_demux_src27_endofpacket),   //           .endofpacket
		.src28_ready         (cmd_xbar_demux_src28_ready),         //      src28.ready
		.src28_valid         (cmd_xbar_demux_src28_valid),         //           .valid
		.src28_data          (cmd_xbar_demux_src28_data),          //           .data
		.src28_channel       (cmd_xbar_demux_src28_channel),       //           .channel
		.src28_startofpacket (cmd_xbar_demux_src28_startofpacket), //           .startofpacket
		.src28_endofpacket   (cmd_xbar_demux_src28_endofpacket),   //           .endofpacket
		.src29_ready         (cmd_xbar_demux_src29_ready),         //      src29.ready
		.src29_valid         (cmd_xbar_demux_src29_valid),         //           .valid
		.src29_data          (cmd_xbar_demux_src29_data),          //           .data
		.src29_channel       (cmd_xbar_demux_src29_channel),       //           .channel
		.src29_startofpacket (cmd_xbar_demux_src29_startofpacket), //           .startofpacket
		.src29_endofpacket   (cmd_xbar_demux_src29_endofpacket),   //           .endofpacket
		.src30_ready         (cmd_xbar_demux_src30_ready),         //      src30.ready
		.src30_valid         (cmd_xbar_demux_src30_valid),         //           .valid
		.src30_data          (cmd_xbar_demux_src30_data),          //           .data
		.src30_channel       (cmd_xbar_demux_src30_channel),       //           .channel
		.src30_startofpacket (cmd_xbar_demux_src30_startofpacket), //           .startofpacket
		.src30_endofpacket   (cmd_xbar_demux_src30_endofpacket),   //           .endofpacket
		.src31_ready         (cmd_xbar_demux_src31_ready),         //      src31.ready
		.src31_valid         (cmd_xbar_demux_src31_valid),         //           .valid
		.src31_data          (cmd_xbar_demux_src31_data),          //           .data
		.src31_channel       (cmd_xbar_demux_src31_channel),       //           .channel
		.src31_startofpacket (cmd_xbar_demux_src31_startofpacket), //           .startofpacket
		.src31_endofpacket   (cmd_xbar_demux_src31_endofpacket),   //           .endofpacket
		.src32_ready         (cmd_xbar_demux_src32_ready),         //      src32.ready
		.src32_valid         (cmd_xbar_demux_src32_valid),         //           .valid
		.src32_data          (cmd_xbar_demux_src32_data),          //           .data
		.src32_channel       (cmd_xbar_demux_src32_channel),       //           .channel
		.src32_startofpacket (cmd_xbar_demux_src32_startofpacket), //           .startofpacket
		.src32_endofpacket   (cmd_xbar_demux_src32_endofpacket),   //           .endofpacket
		.src33_ready         (cmd_xbar_demux_src33_ready),         //      src33.ready
		.src33_valid         (cmd_xbar_demux_src33_valid),         //           .valid
		.src33_data          (cmd_xbar_demux_src33_data),          //           .data
		.src33_channel       (cmd_xbar_demux_src33_channel),       //           .channel
		.src33_startofpacket (cmd_xbar_demux_src33_startofpacket), //           .startofpacket
		.src33_endofpacket   (cmd_xbar_demux_src33_endofpacket),   //           .endofpacket
		.src34_ready         (cmd_xbar_demux_src34_ready),         //      src34.ready
		.src34_valid         (cmd_xbar_demux_src34_valid),         //           .valid
		.src34_data          (cmd_xbar_demux_src34_data),          //           .data
		.src34_channel       (cmd_xbar_demux_src34_channel),       //           .channel
		.src34_startofpacket (cmd_xbar_demux_src34_startofpacket), //           .startofpacket
		.src34_endofpacket   (cmd_xbar_demux_src34_endofpacket),   //           .endofpacket
		.src35_ready         (cmd_xbar_demux_src35_ready),         //      src35.ready
		.src35_valid         (cmd_xbar_demux_src35_valid),         //           .valid
		.src35_data          (cmd_xbar_demux_src35_data),          //           .data
		.src35_channel       (cmd_xbar_demux_src35_channel),       //           .channel
		.src35_startofpacket (cmd_xbar_demux_src35_startofpacket), //           .startofpacket
		.src35_endofpacket   (cmd_xbar_demux_src35_endofpacket),   //           .endofpacket
		.src36_ready         (cmd_xbar_demux_src36_ready),         //      src36.ready
		.src36_valid         (cmd_xbar_demux_src36_valid),         //           .valid
		.src36_data          (cmd_xbar_demux_src36_data),          //           .data
		.src36_channel       (cmd_xbar_demux_src36_channel),       //           .channel
		.src36_startofpacket (cmd_xbar_demux_src36_startofpacket), //           .startofpacket
		.src36_endofpacket   (cmd_xbar_demux_src36_endofpacket),   //           .endofpacket
		.src37_ready         (cmd_xbar_demux_src37_ready),         //      src37.ready
		.src37_valid         (cmd_xbar_demux_src37_valid),         //           .valid
		.src37_data          (cmd_xbar_demux_src37_data),          //           .data
		.src37_channel       (cmd_xbar_demux_src37_channel),       //           .channel
		.src37_startofpacket (cmd_xbar_demux_src37_startofpacket), //           .startofpacket
		.src37_endofpacket   (cmd_xbar_demux_src37_endofpacket),   //           .endofpacket
		.src38_ready         (cmd_xbar_demux_src38_ready),         //      src38.ready
		.src38_valid         (cmd_xbar_demux_src38_valid),         //           .valid
		.src38_data          (cmd_xbar_demux_src38_data),          //           .data
		.src38_channel       (cmd_xbar_demux_src38_channel),       //           .channel
		.src38_startofpacket (cmd_xbar_demux_src38_startofpacket), //           .startofpacket
		.src38_endofpacket   (cmd_xbar_demux_src38_endofpacket),   //           .endofpacket
		.src39_ready         (cmd_xbar_demux_src39_ready),         //      src39.ready
		.src39_valid         (cmd_xbar_demux_src39_valid),         //           .valid
		.src39_data          (cmd_xbar_demux_src39_data),          //           .data
		.src39_channel       (cmd_xbar_demux_src39_channel),       //           .channel
		.src39_startofpacket (cmd_xbar_demux_src39_startofpacket), //           .startofpacket
		.src39_endofpacket   (cmd_xbar_demux_src39_endofpacket),   //           .endofpacket
		.src40_ready         (cmd_xbar_demux_src40_ready),         //      src40.ready
		.src40_valid         (cmd_xbar_demux_src40_valid),         //           .valid
		.src40_data          (cmd_xbar_demux_src40_data),          //           .data
		.src40_channel       (cmd_xbar_demux_src40_channel),       //           .channel
		.src40_startofpacket (cmd_xbar_demux_src40_startofpacket), //           .startofpacket
		.src40_endofpacket   (cmd_xbar_demux_src40_endofpacket),   //           .endofpacket
		.src41_ready         (cmd_xbar_demux_src41_ready),         //      src41.ready
		.src41_valid         (cmd_xbar_demux_src41_valid),         //           .valid
		.src41_data          (cmd_xbar_demux_src41_data),          //           .data
		.src41_channel       (cmd_xbar_demux_src41_channel),       //           .channel
		.src41_startofpacket (cmd_xbar_demux_src41_startofpacket), //           .startofpacket
		.src41_endofpacket   (cmd_xbar_demux_src41_endofpacket),   //           .endofpacket
		.src42_ready         (cmd_xbar_demux_src42_ready),         //      src42.ready
		.src42_valid         (cmd_xbar_demux_src42_valid),         //           .valid
		.src42_data          (cmd_xbar_demux_src42_data),          //           .data
		.src42_channel       (cmd_xbar_demux_src42_channel),       //           .channel
		.src42_startofpacket (cmd_xbar_demux_src42_startofpacket), //           .startofpacket
		.src42_endofpacket   (cmd_xbar_demux_src42_endofpacket),   //           .endofpacket
		.src43_ready         (cmd_xbar_demux_src43_ready),         //      src43.ready
		.src43_valid         (cmd_xbar_demux_src43_valid),         //           .valid
		.src43_data          (cmd_xbar_demux_src43_data),          //           .data
		.src43_channel       (cmd_xbar_demux_src43_channel),       //           .channel
		.src43_startofpacket (cmd_xbar_demux_src43_startofpacket), //           .startofpacket
		.src43_endofpacket   (cmd_xbar_demux_src43_endofpacket),   //           .endofpacket
		.src44_ready         (cmd_xbar_demux_src44_ready),         //      src44.ready
		.src44_valid         (cmd_xbar_demux_src44_valid),         //           .valid
		.src44_data          (cmd_xbar_demux_src44_data),          //           .data
		.src44_channel       (cmd_xbar_demux_src44_channel),       //           .channel
		.src44_startofpacket (cmd_xbar_demux_src44_startofpacket), //           .startofpacket
		.src44_endofpacket   (cmd_xbar_demux_src44_endofpacket),   //           .endofpacket
		.src45_ready         (cmd_xbar_demux_src45_ready),         //      src45.ready
		.src45_valid         (cmd_xbar_demux_src45_valid),         //           .valid
		.src45_data          (cmd_xbar_demux_src45_data),          //           .data
		.src45_channel       (cmd_xbar_demux_src45_channel),       //           .channel
		.src45_startofpacket (cmd_xbar_demux_src45_startofpacket), //           .startofpacket
		.src45_endofpacket   (cmd_xbar_demux_src45_endofpacket),   //           .endofpacket
		.src46_ready         (cmd_xbar_demux_src46_ready),         //      src46.ready
		.src46_valid         (cmd_xbar_demux_src46_valid),         //           .valid
		.src46_data          (cmd_xbar_demux_src46_data),          //           .data
		.src46_channel       (cmd_xbar_demux_src46_channel),       //           .channel
		.src46_startofpacket (cmd_xbar_demux_src46_startofpacket), //           .startofpacket
		.src46_endofpacket   (cmd_xbar_demux_src46_endofpacket),   //           .endofpacket
		.src47_ready         (cmd_xbar_demux_src47_ready),         //      src47.ready
		.src47_valid         (cmd_xbar_demux_src47_valid),         //           .valid
		.src47_data          (cmd_xbar_demux_src47_data),          //           .data
		.src47_channel       (cmd_xbar_demux_src47_channel),       //           .channel
		.src47_startofpacket (cmd_xbar_demux_src47_startofpacket), //           .startofpacket
		.src47_endofpacket   (cmd_xbar_demux_src47_endofpacket),   //           .endofpacket
		.src48_ready         (cmd_xbar_demux_src48_ready),         //      src48.ready
		.src48_valid         (cmd_xbar_demux_src48_valid),         //           .valid
		.src48_data          (cmd_xbar_demux_src48_data),          //           .data
		.src48_channel       (cmd_xbar_demux_src48_channel),       //           .channel
		.src48_startofpacket (cmd_xbar_demux_src48_startofpacket), //           .startofpacket
		.src48_endofpacket   (cmd_xbar_demux_src48_endofpacket),   //           .endofpacket
		.src49_ready         (cmd_xbar_demux_src49_ready),         //      src49.ready
		.src49_valid         (cmd_xbar_demux_src49_valid),         //           .valid
		.src49_data          (cmd_xbar_demux_src49_data),          //           .data
		.src49_channel       (cmd_xbar_demux_src49_channel),       //           .channel
		.src49_startofpacket (cmd_xbar_demux_src49_startofpacket), //           .startofpacket
		.src49_endofpacket   (cmd_xbar_demux_src49_endofpacket),   //           .endofpacket
		.src50_ready         (cmd_xbar_demux_src50_ready),         //      src50.ready
		.src50_valid         (cmd_xbar_demux_src50_valid),         //           .valid
		.src50_data          (cmd_xbar_demux_src50_data),          //           .data
		.src50_channel       (cmd_xbar_demux_src50_channel),       //           .channel
		.src50_startofpacket (cmd_xbar_demux_src50_startofpacket), //           .startofpacket
		.src50_endofpacket   (cmd_xbar_demux_src50_endofpacket),   //           .endofpacket
		.src51_ready         (cmd_xbar_demux_src51_ready),         //      src51.ready
		.src51_valid         (cmd_xbar_demux_src51_valid),         //           .valid
		.src51_data          (cmd_xbar_demux_src51_data),          //           .data
		.src51_channel       (cmd_xbar_demux_src51_channel),       //           .channel
		.src51_startofpacket (cmd_xbar_demux_src51_startofpacket), //           .startofpacket
		.src51_endofpacket   (cmd_xbar_demux_src51_endofpacket),   //           .endofpacket
		.src52_ready         (cmd_xbar_demux_src52_ready),         //      src52.ready
		.src52_valid         (cmd_xbar_demux_src52_valid),         //           .valid
		.src52_data          (cmd_xbar_demux_src52_data),          //           .data
		.src52_channel       (cmd_xbar_demux_src52_channel),       //           .channel
		.src52_startofpacket (cmd_xbar_demux_src52_startofpacket), //           .startofpacket
		.src52_endofpacket   (cmd_xbar_demux_src52_endofpacket),   //           .endofpacket
		.src53_ready         (cmd_xbar_demux_src53_ready),         //      src53.ready
		.src53_valid         (cmd_xbar_demux_src53_valid),         //           .valid
		.src53_data          (cmd_xbar_demux_src53_data),          //           .data
		.src53_channel       (cmd_xbar_demux_src53_channel),       //           .channel
		.src53_startofpacket (cmd_xbar_demux_src53_startofpacket), //           .startofpacket
		.src53_endofpacket   (cmd_xbar_demux_src53_endofpacket),   //           .endofpacket
		.src54_ready         (cmd_xbar_demux_src54_ready),         //      src54.ready
		.src54_valid         (cmd_xbar_demux_src54_valid),         //           .valid
		.src54_data          (cmd_xbar_demux_src54_data),          //           .data
		.src54_channel       (cmd_xbar_demux_src54_channel),       //           .channel
		.src54_startofpacket (cmd_xbar_demux_src54_startofpacket), //           .startofpacket
		.src54_endofpacket   (cmd_xbar_demux_src54_endofpacket),   //           .endofpacket
		.src55_ready         (cmd_xbar_demux_src55_ready),         //      src55.ready
		.src55_valid         (cmd_xbar_demux_src55_valid),         //           .valid
		.src55_data          (cmd_xbar_demux_src55_data),          //           .data
		.src55_channel       (cmd_xbar_demux_src55_channel),       //           .channel
		.src55_startofpacket (cmd_xbar_demux_src55_startofpacket), //           .startofpacket
		.src55_endofpacket   (cmd_xbar_demux_src55_endofpacket),   //           .endofpacket
		.src56_ready         (cmd_xbar_demux_src56_ready),         //      src56.ready
		.src56_valid         (cmd_xbar_demux_src56_valid),         //           .valid
		.src56_data          (cmd_xbar_demux_src56_data),          //           .data
		.src56_channel       (cmd_xbar_demux_src56_channel),       //           .channel
		.src56_startofpacket (cmd_xbar_demux_src56_startofpacket), //           .startofpacket
		.src56_endofpacket   (cmd_xbar_demux_src56_endofpacket),   //           .endofpacket
		.src57_ready         (cmd_xbar_demux_src57_ready),         //      src57.ready
		.src57_valid         (cmd_xbar_demux_src57_valid),         //           .valid
		.src57_data          (cmd_xbar_demux_src57_data),          //           .data
		.src57_channel       (cmd_xbar_demux_src57_channel),       //           .channel
		.src57_startofpacket (cmd_xbar_demux_src57_startofpacket), //           .startofpacket
		.src57_endofpacket   (cmd_xbar_demux_src57_endofpacket)    //           .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux (
		.clk                (sam9_mclk_clk),                     //       clk.clk
		.reset              (sam9_mrst_reset),                   // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_007 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_008 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_005_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_005_src_channel),         //          .channel
		.sink_data          (width_adapter_005_src_data),            //          .data
		.sink_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_005_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_009 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_007_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_007_src_channel),         //          .channel
		.sink_data          (width_adapter_007_src_data),            //          .data
		.sink_startofpacket (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_007_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_010 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_009_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_009_src_channel),         //          .channel
		.sink_data          (width_adapter_009_src_data),            //          .data
		.sink_startofpacket (width_adapter_009_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_009_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_009_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_011 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_011_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_011_src_channel),         //          .channel
		.sink_data          (width_adapter_011_src_data),            //          .data
		.sink_startofpacket (width_adapter_011_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_011_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_011_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_012 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_013_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_013_src_channel),         //          .channel
		.sink_data          (width_adapter_013_src_data),            //          .data
		.sink_startofpacket (width_adapter_013_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_013_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_013_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_013 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_015_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_015_src_channel),         //          .channel
		.sink_data          (width_adapter_015_src_data),            //          .data
		.sink_startofpacket (width_adapter_015_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_015_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_015_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_014 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_017_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_017_src_channel),         //          .channel
		.sink_data          (width_adapter_017_src_data),            //          .data
		.sink_startofpacket (width_adapter_017_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_017_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_017_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_015 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_019_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_019_src_channel),         //          .channel
		.sink_data          (width_adapter_019_src_data),            //          .data
		.sink_startofpacket (width_adapter_019_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_019_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_019_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_016 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_021_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_021_src_channel),         //          .channel
		.sink_data          (width_adapter_021_src_data),            //          .data
		.sink_startofpacket (width_adapter_021_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_021_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_021_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_017 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_023_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_023_src_channel),         //          .channel
		.sink_data          (width_adapter_023_src_data),            //          .data
		.sink_startofpacket (width_adapter_023_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_023_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_023_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_018 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_025_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_025_src_channel),         //          .channel
		.sink_data          (width_adapter_025_src_data),            //          .data
		.sink_startofpacket (width_adapter_025_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_025_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_025_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_019 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_027_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_027_src_channel),         //          .channel
		.sink_data          (width_adapter_027_src_data),            //          .data
		.sink_startofpacket (width_adapter_027_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_027_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_027_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_020 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_029_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_029_src_channel),         //          .channel
		.sink_data          (width_adapter_029_src_data),            //          .data
		.sink_startofpacket (width_adapter_029_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_029_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_029_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_021 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_031_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_031_src_channel),         //          .channel
		.sink_data          (width_adapter_031_src_data),            //          .data
		.sink_startofpacket (width_adapter_031_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_031_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_031_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_022 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_033_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_033_src_channel),         //          .channel
		.sink_data          (width_adapter_033_src_data),            //          .data
		.sink_startofpacket (width_adapter_033_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_033_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_033_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_023 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_035_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_035_src_channel),         //          .channel
		.sink_data          (width_adapter_035_src_data),            //          .data
		.sink_startofpacket (width_adapter_035_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_035_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_035_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_024 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_037_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_037_src_channel),         //          .channel
		.sink_data          (width_adapter_037_src_data),            //          .data
		.sink_startofpacket (width_adapter_037_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_037_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_037_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_025 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_039_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_039_src_channel),         //          .channel
		.sink_data          (width_adapter_039_src_data),            //          .data
		.sink_startofpacket (width_adapter_039_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_039_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_039_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_026 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_041_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_041_src_channel),         //          .channel
		.sink_data          (width_adapter_041_src_data),            //          .data
		.sink_startofpacket (width_adapter_041_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_041_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_041_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_026_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_026_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_027 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_043_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_043_src_channel),         //          .channel
		.sink_data          (width_adapter_043_src_data),            //          .data
		.sink_startofpacket (width_adapter_043_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_043_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_043_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_027_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_027_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_028 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_045_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_045_src_channel),         //          .channel
		.sink_data          (width_adapter_045_src_data),            //          .data
		.sink_startofpacket (width_adapter_045_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_045_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_045_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_028_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_029 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_047_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_047_src_channel),         //          .channel
		.sink_data          (width_adapter_047_src_data),            //          .data
		.sink_startofpacket (width_adapter_047_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_047_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_047_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_029_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_030 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_049_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_049_src_channel),         //          .channel
		.sink_data          (width_adapter_049_src_data),            //          .data
		.sink_startofpacket (width_adapter_049_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_049_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_049_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_030_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_030_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_031 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_051_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_051_src_channel),         //          .channel
		.sink_data          (width_adapter_051_src_data),            //          .data
		.sink_startofpacket (width_adapter_051_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_051_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_051_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_031_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_031_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_032 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_053_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_053_src_channel),         //          .channel
		.sink_data          (width_adapter_053_src_data),            //          .data
		.sink_startofpacket (width_adapter_053_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_053_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_053_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_032_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_032_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_033 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_055_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_055_src_channel),         //          .channel
		.sink_data          (width_adapter_055_src_data),            //          .data
		.sink_startofpacket (width_adapter_055_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_055_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_055_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_033_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_033_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_034 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_057_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_057_src_channel),         //          .channel
		.sink_data          (width_adapter_057_src_data),            //          .data
		.sink_startofpacket (width_adapter_057_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_057_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_057_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_034_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_034_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_035 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_059_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_059_src_channel),         //          .channel
		.sink_data          (width_adapter_059_src_data),            //          .data
		.sink_startofpacket (width_adapter_059_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_059_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_059_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_035_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_035_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_036 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_061_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_061_src_channel),         //          .channel
		.sink_data          (width_adapter_061_src_data),            //          .data
		.sink_startofpacket (width_adapter_061_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_061_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_061_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_036_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_036_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_037 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_063_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_063_src_channel),         //          .channel
		.sink_data          (width_adapter_063_src_data),            //          .data
		.sink_startofpacket (width_adapter_063_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_063_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_063_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_037_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_037_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_037_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_037_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_037_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_038 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_065_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_065_src_channel),         //          .channel
		.sink_data          (width_adapter_065_src_data),            //          .data
		.sink_startofpacket (width_adapter_065_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_065_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_065_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_038_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_038_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_038_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_038_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_038_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_038_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_039 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_067_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_067_src_channel),         //          .channel
		.sink_data          (width_adapter_067_src_data),            //          .data
		.sink_startofpacket (width_adapter_067_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_067_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_067_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_039_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_039_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_039_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_039_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_039_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_039_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_040 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_069_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_069_src_channel),         //          .channel
		.sink_data          (width_adapter_069_src_data),            //          .data
		.sink_startofpacket (width_adapter_069_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_069_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_069_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_040_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_040_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_040_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_040_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_040_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_040_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_041 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_071_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_071_src_channel),         //          .channel
		.sink_data          (width_adapter_071_src_data),            //          .data
		.sink_startofpacket (width_adapter_071_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_071_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_071_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_041_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_041_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_041_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_041_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_041_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_041_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_042 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_073_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_073_src_channel),         //          .channel
		.sink_data          (width_adapter_073_src_data),            //          .data
		.sink_startofpacket (width_adapter_073_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_073_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_073_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_042_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_042_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_042_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_042_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_042_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_042_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_043 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_075_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_075_src_channel),         //          .channel
		.sink_data          (width_adapter_075_src_data),            //          .data
		.sink_startofpacket (width_adapter_075_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_075_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_075_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_043_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_043_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_043_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_043_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_043_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_043_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_044 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_077_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_077_src_channel),         //          .channel
		.sink_data          (width_adapter_077_src_data),            //          .data
		.sink_startofpacket (width_adapter_077_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_077_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_077_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_044_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_044_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_044_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_044_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_044_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_044_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_045 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_079_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_079_src_channel),         //          .channel
		.sink_data          (width_adapter_079_src_data),            //          .data
		.sink_startofpacket (width_adapter_079_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_079_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_079_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_045_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_045_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_045_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_045_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_045_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_045_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_046 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_081_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_081_src_channel),         //          .channel
		.sink_data          (width_adapter_081_src_data),            //          .data
		.sink_startofpacket (width_adapter_081_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_081_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_081_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_046_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_046_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_046_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_046_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_046_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_046_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_047 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_083_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_083_src_channel),         //          .channel
		.sink_data          (width_adapter_083_src_data),            //          .data
		.sink_startofpacket (width_adapter_083_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_083_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_083_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_047_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_047_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_047_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_047_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_047_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_047_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_048 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_085_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_085_src_channel),         //          .channel
		.sink_data          (width_adapter_085_src_data),            //          .data
		.sink_startofpacket (width_adapter_085_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_085_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_085_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_048_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_048_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_048_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_048_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_048_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_048_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_049 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_087_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_087_src_channel),         //          .channel
		.sink_data          (width_adapter_087_src_data),            //          .data
		.sink_startofpacket (width_adapter_087_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_087_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_087_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_049_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_049_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_049_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_049_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_049_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_049_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_050 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_089_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_089_src_channel),         //          .channel
		.sink_data          (width_adapter_089_src_data),            //          .data
		.sink_startofpacket (width_adapter_089_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_089_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_089_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_050_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_050_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_050_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_050_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_050_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_050_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_051 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_091_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_091_src_channel),         //          .channel
		.sink_data          (width_adapter_091_src_data),            //          .data
		.sink_startofpacket (width_adapter_091_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_091_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_091_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_051_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_051_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_051_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_051_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_051_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_051_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_052 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_093_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_093_src_channel),         //          .channel
		.sink_data          (width_adapter_093_src_data),            //          .data
		.sink_startofpacket (width_adapter_093_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_093_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_093_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_052_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_052_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_052_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_052_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_052_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_052_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_053 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_095_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_095_src_channel),         //          .channel
		.sink_data          (width_adapter_095_src_data),            //          .data
		.sink_startofpacket (width_adapter_095_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_095_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_095_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_053_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_053_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_053_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_053_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_053_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_053_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_054 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_097_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_097_src_channel),         //          .channel
		.sink_data          (width_adapter_097_src_data),            //          .data
		.sink_startofpacket (width_adapter_097_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_097_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_097_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_054_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_054_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_054_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_054_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_054_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_054_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_055 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_099_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_099_src_channel),         //          .channel
		.sink_data          (width_adapter_099_src_data),            //          .data
		.sink_startofpacket (width_adapter_099_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_099_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_099_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_055_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_055_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_055_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_055_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_055_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_055_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_056 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_101_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_101_src_channel),         //          .channel
		.sink_data          (width_adapter_101_src_data),            //          .data
		.sink_startofpacket (width_adapter_101_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_101_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_101_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_056_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_056_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_056_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_056_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_056_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_056_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_057 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (width_adapter_103_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_103_src_channel),         //          .channel
		.sink_data          (width_adapter_103_src_data),            //          .data
		.sink_startofpacket (width_adapter_103_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_103_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_103_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_057_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_057_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_057_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_057_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_057_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_057_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_mux rsp_xbar_mux (
		.clk                  (sam9_mclk_clk),                         //       clk.clk
		.reset                (sam9_mrst_reset),                       // clk_reset.reset
		.src_ready            (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid            (rsp_xbar_mux_src_valid),                //          .valid
		.src_data             (rsp_xbar_mux_src_data),                 //          .data
		.src_channel          (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket    (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_021_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_022_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink23_ready         (rsp_xbar_demux_023_src0_ready),         //    sink23.ready
		.sink23_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink23_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink23_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink23_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink23_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink24_ready         (rsp_xbar_demux_024_src0_ready),         //    sink24.ready
		.sink24_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink24_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink24_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink24_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink24_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink25_ready         (rsp_xbar_demux_025_src0_ready),         //    sink25.ready
		.sink25_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.sink25_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.sink25_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.sink25_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.sink25_endofpacket   (rsp_xbar_demux_025_src0_endofpacket),   //          .endofpacket
		.sink26_ready         (rsp_xbar_demux_026_src0_ready),         //    sink26.ready
		.sink26_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.sink26_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.sink26_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.sink26_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.sink26_endofpacket   (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.sink27_ready         (rsp_xbar_demux_027_src0_ready),         //    sink27.ready
		.sink27_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.sink27_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.sink27_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.sink27_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.sink27_endofpacket   (rsp_xbar_demux_027_src0_endofpacket),   //          .endofpacket
		.sink28_ready         (rsp_xbar_demux_028_src0_ready),         //    sink28.ready
		.sink28_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.sink28_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.sink28_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.sink28_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.sink28_endofpacket   (rsp_xbar_demux_028_src0_endofpacket),   //          .endofpacket
		.sink29_ready         (rsp_xbar_demux_029_src0_ready),         //    sink29.ready
		.sink29_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.sink29_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.sink29_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.sink29_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.sink29_endofpacket   (rsp_xbar_demux_029_src0_endofpacket),   //          .endofpacket
		.sink30_ready         (rsp_xbar_demux_030_src0_ready),         //    sink30.ready
		.sink30_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.sink30_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.sink30_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.sink30_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.sink30_endofpacket   (rsp_xbar_demux_030_src0_endofpacket),   //          .endofpacket
		.sink31_ready         (rsp_xbar_demux_031_src0_ready),         //    sink31.ready
		.sink31_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.sink31_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.sink31_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.sink31_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.sink31_endofpacket   (rsp_xbar_demux_031_src0_endofpacket),   //          .endofpacket
		.sink32_ready         (rsp_xbar_demux_032_src0_ready),         //    sink32.ready
		.sink32_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.sink32_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.sink32_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.sink32_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.sink32_endofpacket   (rsp_xbar_demux_032_src0_endofpacket),   //          .endofpacket
		.sink33_ready         (rsp_xbar_demux_033_src0_ready),         //    sink33.ready
		.sink33_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.sink33_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.sink33_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.sink33_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.sink33_endofpacket   (rsp_xbar_demux_033_src0_endofpacket),   //          .endofpacket
		.sink34_ready         (rsp_xbar_demux_034_src0_ready),         //    sink34.ready
		.sink34_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.sink34_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.sink34_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.sink34_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.sink34_endofpacket   (rsp_xbar_demux_034_src0_endofpacket),   //          .endofpacket
		.sink35_ready         (rsp_xbar_demux_035_src0_ready),         //    sink35.ready
		.sink35_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.sink35_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.sink35_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.sink35_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.sink35_endofpacket   (rsp_xbar_demux_035_src0_endofpacket),   //          .endofpacket
		.sink36_ready         (rsp_xbar_demux_036_src0_ready),         //    sink36.ready
		.sink36_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.sink36_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.sink36_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.sink36_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.sink36_endofpacket   (rsp_xbar_demux_036_src0_endofpacket),   //          .endofpacket
		.sink37_ready         (rsp_xbar_demux_037_src0_ready),         //    sink37.ready
		.sink37_valid         (rsp_xbar_demux_037_src0_valid),         //          .valid
		.sink37_channel       (rsp_xbar_demux_037_src0_channel),       //          .channel
		.sink37_data          (rsp_xbar_demux_037_src0_data),          //          .data
		.sink37_startofpacket (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.sink37_endofpacket   (rsp_xbar_demux_037_src0_endofpacket),   //          .endofpacket
		.sink38_ready         (rsp_xbar_demux_038_src0_ready),         //    sink38.ready
		.sink38_valid         (rsp_xbar_demux_038_src0_valid),         //          .valid
		.sink38_channel       (rsp_xbar_demux_038_src0_channel),       //          .channel
		.sink38_data          (rsp_xbar_demux_038_src0_data),          //          .data
		.sink38_startofpacket (rsp_xbar_demux_038_src0_startofpacket), //          .startofpacket
		.sink38_endofpacket   (rsp_xbar_demux_038_src0_endofpacket),   //          .endofpacket
		.sink39_ready         (rsp_xbar_demux_039_src0_ready),         //    sink39.ready
		.sink39_valid         (rsp_xbar_demux_039_src0_valid),         //          .valid
		.sink39_channel       (rsp_xbar_demux_039_src0_channel),       //          .channel
		.sink39_data          (rsp_xbar_demux_039_src0_data),          //          .data
		.sink39_startofpacket (rsp_xbar_demux_039_src0_startofpacket), //          .startofpacket
		.sink39_endofpacket   (rsp_xbar_demux_039_src0_endofpacket),   //          .endofpacket
		.sink40_ready         (rsp_xbar_demux_040_src0_ready),         //    sink40.ready
		.sink40_valid         (rsp_xbar_demux_040_src0_valid),         //          .valid
		.sink40_channel       (rsp_xbar_demux_040_src0_channel),       //          .channel
		.sink40_data          (rsp_xbar_demux_040_src0_data),          //          .data
		.sink40_startofpacket (rsp_xbar_demux_040_src0_startofpacket), //          .startofpacket
		.sink40_endofpacket   (rsp_xbar_demux_040_src0_endofpacket),   //          .endofpacket
		.sink41_ready         (rsp_xbar_demux_041_src0_ready),         //    sink41.ready
		.sink41_valid         (rsp_xbar_demux_041_src0_valid),         //          .valid
		.sink41_channel       (rsp_xbar_demux_041_src0_channel),       //          .channel
		.sink41_data          (rsp_xbar_demux_041_src0_data),          //          .data
		.sink41_startofpacket (rsp_xbar_demux_041_src0_startofpacket), //          .startofpacket
		.sink41_endofpacket   (rsp_xbar_demux_041_src0_endofpacket),   //          .endofpacket
		.sink42_ready         (rsp_xbar_demux_042_src0_ready),         //    sink42.ready
		.sink42_valid         (rsp_xbar_demux_042_src0_valid),         //          .valid
		.sink42_channel       (rsp_xbar_demux_042_src0_channel),       //          .channel
		.sink42_data          (rsp_xbar_demux_042_src0_data),          //          .data
		.sink42_startofpacket (rsp_xbar_demux_042_src0_startofpacket), //          .startofpacket
		.sink42_endofpacket   (rsp_xbar_demux_042_src0_endofpacket),   //          .endofpacket
		.sink43_ready         (rsp_xbar_demux_043_src0_ready),         //    sink43.ready
		.sink43_valid         (rsp_xbar_demux_043_src0_valid),         //          .valid
		.sink43_channel       (rsp_xbar_demux_043_src0_channel),       //          .channel
		.sink43_data          (rsp_xbar_demux_043_src0_data),          //          .data
		.sink43_startofpacket (rsp_xbar_demux_043_src0_startofpacket), //          .startofpacket
		.sink43_endofpacket   (rsp_xbar_demux_043_src0_endofpacket),   //          .endofpacket
		.sink44_ready         (rsp_xbar_demux_044_src0_ready),         //    sink44.ready
		.sink44_valid         (rsp_xbar_demux_044_src0_valid),         //          .valid
		.sink44_channel       (rsp_xbar_demux_044_src0_channel),       //          .channel
		.sink44_data          (rsp_xbar_demux_044_src0_data),          //          .data
		.sink44_startofpacket (rsp_xbar_demux_044_src0_startofpacket), //          .startofpacket
		.sink44_endofpacket   (rsp_xbar_demux_044_src0_endofpacket),   //          .endofpacket
		.sink45_ready         (rsp_xbar_demux_045_src0_ready),         //    sink45.ready
		.sink45_valid         (rsp_xbar_demux_045_src0_valid),         //          .valid
		.sink45_channel       (rsp_xbar_demux_045_src0_channel),       //          .channel
		.sink45_data          (rsp_xbar_demux_045_src0_data),          //          .data
		.sink45_startofpacket (rsp_xbar_demux_045_src0_startofpacket), //          .startofpacket
		.sink45_endofpacket   (rsp_xbar_demux_045_src0_endofpacket),   //          .endofpacket
		.sink46_ready         (rsp_xbar_demux_046_src0_ready),         //    sink46.ready
		.sink46_valid         (rsp_xbar_demux_046_src0_valid),         //          .valid
		.sink46_channel       (rsp_xbar_demux_046_src0_channel),       //          .channel
		.sink46_data          (rsp_xbar_demux_046_src0_data),          //          .data
		.sink46_startofpacket (rsp_xbar_demux_046_src0_startofpacket), //          .startofpacket
		.sink46_endofpacket   (rsp_xbar_demux_046_src0_endofpacket),   //          .endofpacket
		.sink47_ready         (rsp_xbar_demux_047_src0_ready),         //    sink47.ready
		.sink47_valid         (rsp_xbar_demux_047_src0_valid),         //          .valid
		.sink47_channel       (rsp_xbar_demux_047_src0_channel),       //          .channel
		.sink47_data          (rsp_xbar_demux_047_src0_data),          //          .data
		.sink47_startofpacket (rsp_xbar_demux_047_src0_startofpacket), //          .startofpacket
		.sink47_endofpacket   (rsp_xbar_demux_047_src0_endofpacket),   //          .endofpacket
		.sink48_ready         (rsp_xbar_demux_048_src0_ready),         //    sink48.ready
		.sink48_valid         (rsp_xbar_demux_048_src0_valid),         //          .valid
		.sink48_channel       (rsp_xbar_demux_048_src0_channel),       //          .channel
		.sink48_data          (rsp_xbar_demux_048_src0_data),          //          .data
		.sink48_startofpacket (rsp_xbar_demux_048_src0_startofpacket), //          .startofpacket
		.sink48_endofpacket   (rsp_xbar_demux_048_src0_endofpacket),   //          .endofpacket
		.sink49_ready         (rsp_xbar_demux_049_src0_ready),         //    sink49.ready
		.sink49_valid         (rsp_xbar_demux_049_src0_valid),         //          .valid
		.sink49_channel       (rsp_xbar_demux_049_src0_channel),       //          .channel
		.sink49_data          (rsp_xbar_demux_049_src0_data),          //          .data
		.sink49_startofpacket (rsp_xbar_demux_049_src0_startofpacket), //          .startofpacket
		.sink49_endofpacket   (rsp_xbar_demux_049_src0_endofpacket),   //          .endofpacket
		.sink50_ready         (rsp_xbar_demux_050_src0_ready),         //    sink50.ready
		.sink50_valid         (rsp_xbar_demux_050_src0_valid),         //          .valid
		.sink50_channel       (rsp_xbar_demux_050_src0_channel),       //          .channel
		.sink50_data          (rsp_xbar_demux_050_src0_data),          //          .data
		.sink50_startofpacket (rsp_xbar_demux_050_src0_startofpacket), //          .startofpacket
		.sink50_endofpacket   (rsp_xbar_demux_050_src0_endofpacket),   //          .endofpacket
		.sink51_ready         (rsp_xbar_demux_051_src0_ready),         //    sink51.ready
		.sink51_valid         (rsp_xbar_demux_051_src0_valid),         //          .valid
		.sink51_channel       (rsp_xbar_demux_051_src0_channel),       //          .channel
		.sink51_data          (rsp_xbar_demux_051_src0_data),          //          .data
		.sink51_startofpacket (rsp_xbar_demux_051_src0_startofpacket), //          .startofpacket
		.sink51_endofpacket   (rsp_xbar_demux_051_src0_endofpacket),   //          .endofpacket
		.sink52_ready         (rsp_xbar_demux_052_src0_ready),         //    sink52.ready
		.sink52_valid         (rsp_xbar_demux_052_src0_valid),         //          .valid
		.sink52_channel       (rsp_xbar_demux_052_src0_channel),       //          .channel
		.sink52_data          (rsp_xbar_demux_052_src0_data),          //          .data
		.sink52_startofpacket (rsp_xbar_demux_052_src0_startofpacket), //          .startofpacket
		.sink52_endofpacket   (rsp_xbar_demux_052_src0_endofpacket),   //          .endofpacket
		.sink53_ready         (rsp_xbar_demux_053_src0_ready),         //    sink53.ready
		.sink53_valid         (rsp_xbar_demux_053_src0_valid),         //          .valid
		.sink53_channel       (rsp_xbar_demux_053_src0_channel),       //          .channel
		.sink53_data          (rsp_xbar_demux_053_src0_data),          //          .data
		.sink53_startofpacket (rsp_xbar_demux_053_src0_startofpacket), //          .startofpacket
		.sink53_endofpacket   (rsp_xbar_demux_053_src0_endofpacket),   //          .endofpacket
		.sink54_ready         (rsp_xbar_demux_054_src0_ready),         //    sink54.ready
		.sink54_valid         (rsp_xbar_demux_054_src0_valid),         //          .valid
		.sink54_channel       (rsp_xbar_demux_054_src0_channel),       //          .channel
		.sink54_data          (rsp_xbar_demux_054_src0_data),          //          .data
		.sink54_startofpacket (rsp_xbar_demux_054_src0_startofpacket), //          .startofpacket
		.sink54_endofpacket   (rsp_xbar_demux_054_src0_endofpacket),   //          .endofpacket
		.sink55_ready         (rsp_xbar_demux_055_src0_ready),         //    sink55.ready
		.sink55_valid         (rsp_xbar_demux_055_src0_valid),         //          .valid
		.sink55_channel       (rsp_xbar_demux_055_src0_channel),       //          .channel
		.sink55_data          (rsp_xbar_demux_055_src0_data),          //          .data
		.sink55_startofpacket (rsp_xbar_demux_055_src0_startofpacket), //          .startofpacket
		.sink55_endofpacket   (rsp_xbar_demux_055_src0_endofpacket),   //          .endofpacket
		.sink56_ready         (rsp_xbar_demux_056_src0_ready),         //    sink56.ready
		.sink56_valid         (rsp_xbar_demux_056_src0_valid),         //          .valid
		.sink56_channel       (rsp_xbar_demux_056_src0_channel),       //          .channel
		.sink56_data          (rsp_xbar_demux_056_src0_data),          //          .data
		.sink56_startofpacket (rsp_xbar_demux_056_src0_startofpacket), //          .startofpacket
		.sink56_endofpacket   (rsp_xbar_demux_056_src0_endofpacket),   //          .endofpacket
		.sink57_ready         (rsp_xbar_demux_057_src0_ready),         //    sink57.ready
		.sink57_valid         (rsp_xbar_demux_057_src0_valid),         //          .valid
		.sink57_channel       (rsp_xbar_demux_057_src0_channel),       //          .channel
		.sink57_data          (rsp_xbar_demux_057_src0_data),          //          .data
		.sink57_startofpacket (rsp_xbar_demux_057_src0_startofpacket), //          .startofpacket
		.sink57_endofpacket   (rsp_xbar_demux_057_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk               (sam9_mclk_clk),                     //       clk.clk
		.reset             (sam9_mrst_reset),                   // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src6_valid),         //      sink.valid
		.in_channel        (cmd_xbar_demux_src6_channel),       //          .channel
		.in_startofpacket  (cmd_xbar_demux_src6_startofpacket), //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src6_endofpacket),   //          .endofpacket
		.in_ready          (cmd_xbar_demux_src6_ready),         //          .ready
		.in_data           (cmd_xbar_demux_src6_data),          //          .data
		.out_endofpacket   (width_adapter_src_endofpacket),     //       src.endofpacket
		.out_data          (width_adapter_src_data),            //          .data
		.out_channel       (width_adapter_src_channel),         //          .channel
		.out_valid         (width_adapter_src_valid),           //          .valid
		.out_ready         (width_adapter_src_ready),           //          .ready
		.out_startofpacket (width_adapter_src_startofpacket)    //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_006_src_valid),             //      sink.valid
		.in_channel        (id_router_006_src_channel),           //          .channel
		.in_startofpacket  (id_router_006_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_006_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_006_src_ready),             //          .ready
		.in_data           (id_router_006_src_data),              //          .data
		.out_endofpacket   (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_001_src_data),          //          .data
		.out_channel       (width_adapter_001_src_channel),       //          .channel
		.out_valid         (width_adapter_001_src_valid),         //          .valid
		.out_ready         (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket (width_adapter_001_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src7_valid),           //      sink.valid
		.in_channel        (cmd_xbar_demux_src7_channel),         //          .channel
		.in_startofpacket  (cmd_xbar_demux_src7_startofpacket),   //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src7_endofpacket),     //          .endofpacket
		.in_ready          (cmd_xbar_demux_src7_ready),           //          .ready
		.in_data           (cmd_xbar_demux_src7_data),            //          .data
		.out_endofpacket   (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_002_src_data),          //          .data
		.out_channel       (width_adapter_002_src_channel),       //          .channel
		.out_valid         (width_adapter_002_src_valid),         //          .valid
		.out_ready         (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket (width_adapter_002_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_003 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_007_src_valid),             //      sink.valid
		.in_channel        (id_router_007_src_channel),           //          .channel
		.in_startofpacket  (id_router_007_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_007_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_007_src_ready),             //          .ready
		.in_data           (id_router_007_src_data),              //          .data
		.out_endofpacket   (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_003_src_data),          //          .data
		.out_channel       (width_adapter_003_src_channel),       //          .channel
		.out_valid         (width_adapter_003_src_valid),         //          .valid
		.out_ready         (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket (width_adapter_003_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_004 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src8_valid),           //      sink.valid
		.in_channel        (cmd_xbar_demux_src8_channel),         //          .channel
		.in_startofpacket  (cmd_xbar_demux_src8_startofpacket),   //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src8_endofpacket),     //          .endofpacket
		.in_ready          (cmd_xbar_demux_src8_ready),           //          .ready
		.in_data           (cmd_xbar_demux_src8_data),            //          .data
		.out_endofpacket   (width_adapter_004_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_004_src_data),          //          .data
		.out_channel       (width_adapter_004_src_channel),       //          .channel
		.out_valid         (width_adapter_004_src_valid),         //          .valid
		.out_ready         (width_adapter_004_src_ready),         //          .ready
		.out_startofpacket (width_adapter_004_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_005 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_008_src_valid),             //      sink.valid
		.in_channel        (id_router_008_src_channel),           //          .channel
		.in_startofpacket  (id_router_008_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_008_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_008_src_ready),             //          .ready
		.in_data           (id_router_008_src_data),              //          .data
		.out_endofpacket   (width_adapter_005_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_005_src_data),          //          .data
		.out_channel       (width_adapter_005_src_channel),       //          .channel
		.out_valid         (width_adapter_005_src_valid),         //          .valid
		.out_ready         (width_adapter_005_src_ready),         //          .ready
		.out_startofpacket (width_adapter_005_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_006 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src9_valid),           //      sink.valid
		.in_channel        (cmd_xbar_demux_src9_channel),         //          .channel
		.in_startofpacket  (cmd_xbar_demux_src9_startofpacket),   //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src9_endofpacket),     //          .endofpacket
		.in_ready          (cmd_xbar_demux_src9_ready),           //          .ready
		.in_data           (cmd_xbar_demux_src9_data),            //          .data
		.out_endofpacket   (width_adapter_006_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_006_src_data),          //          .data
		.out_channel       (width_adapter_006_src_channel),       //          .channel
		.out_valid         (width_adapter_006_src_valid),         //          .valid
		.out_ready         (width_adapter_006_src_ready),         //          .ready
		.out_startofpacket (width_adapter_006_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_007 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_009_src_valid),             //      sink.valid
		.in_channel        (id_router_009_src_channel),           //          .channel
		.in_startofpacket  (id_router_009_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_009_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_009_src_ready),             //          .ready
		.in_data           (id_router_009_src_data),              //          .data
		.out_endofpacket   (width_adapter_007_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_007_src_data),          //          .data
		.out_channel       (width_adapter_007_src_channel),       //          .channel
		.out_valid         (width_adapter_007_src_valid),         //          .valid
		.out_ready         (width_adapter_007_src_ready),         //          .ready
		.out_startofpacket (width_adapter_007_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_008 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src10_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src10_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src10_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src10_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src10_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src10_data),           //          .data
		.out_endofpacket   (width_adapter_008_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_008_src_data),          //          .data
		.out_channel       (width_adapter_008_src_channel),       //          .channel
		.out_valid         (width_adapter_008_src_valid),         //          .valid
		.out_ready         (width_adapter_008_src_ready),         //          .ready
		.out_startofpacket (width_adapter_008_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_009 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_010_src_valid),             //      sink.valid
		.in_channel        (id_router_010_src_channel),           //          .channel
		.in_startofpacket  (id_router_010_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_010_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_010_src_ready),             //          .ready
		.in_data           (id_router_010_src_data),              //          .data
		.out_endofpacket   (width_adapter_009_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_009_src_data),          //          .data
		.out_channel       (width_adapter_009_src_channel),       //          .channel
		.out_valid         (width_adapter_009_src_valid),         //          .valid
		.out_ready         (width_adapter_009_src_ready),         //          .ready
		.out_startofpacket (width_adapter_009_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_010 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src11_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src11_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src11_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src11_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src11_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src11_data),           //          .data
		.out_endofpacket   (width_adapter_010_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_010_src_data),          //          .data
		.out_channel       (width_adapter_010_src_channel),       //          .channel
		.out_valid         (width_adapter_010_src_valid),         //          .valid
		.out_ready         (width_adapter_010_src_ready),         //          .ready
		.out_startofpacket (width_adapter_010_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_011 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_011_src_valid),             //      sink.valid
		.in_channel        (id_router_011_src_channel),           //          .channel
		.in_startofpacket  (id_router_011_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_011_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_011_src_ready),             //          .ready
		.in_data           (id_router_011_src_data),              //          .data
		.out_endofpacket   (width_adapter_011_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_011_src_data),          //          .data
		.out_channel       (width_adapter_011_src_channel),       //          .channel
		.out_valid         (width_adapter_011_src_valid),         //          .valid
		.out_ready         (width_adapter_011_src_ready),         //          .ready
		.out_startofpacket (width_adapter_011_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_012 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src12_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src12_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src12_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src12_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src12_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src12_data),           //          .data
		.out_endofpacket   (width_adapter_012_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_012_src_data),          //          .data
		.out_channel       (width_adapter_012_src_channel),       //          .channel
		.out_valid         (width_adapter_012_src_valid),         //          .valid
		.out_ready         (width_adapter_012_src_ready),         //          .ready
		.out_startofpacket (width_adapter_012_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_013 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_012_src_valid),             //      sink.valid
		.in_channel        (id_router_012_src_channel),           //          .channel
		.in_startofpacket  (id_router_012_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_012_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_012_src_ready),             //          .ready
		.in_data           (id_router_012_src_data),              //          .data
		.out_endofpacket   (width_adapter_013_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_013_src_data),          //          .data
		.out_channel       (width_adapter_013_src_channel),       //          .channel
		.out_valid         (width_adapter_013_src_valid),         //          .valid
		.out_ready         (width_adapter_013_src_ready),         //          .ready
		.out_startofpacket (width_adapter_013_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_014 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src13_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src13_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src13_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src13_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src13_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src13_data),           //          .data
		.out_endofpacket   (width_adapter_014_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_014_src_data),          //          .data
		.out_channel       (width_adapter_014_src_channel),       //          .channel
		.out_valid         (width_adapter_014_src_valid),         //          .valid
		.out_ready         (width_adapter_014_src_ready),         //          .ready
		.out_startofpacket (width_adapter_014_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_015 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_013_src_valid),             //      sink.valid
		.in_channel        (id_router_013_src_channel),           //          .channel
		.in_startofpacket  (id_router_013_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_013_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_013_src_ready),             //          .ready
		.in_data           (id_router_013_src_data),              //          .data
		.out_endofpacket   (width_adapter_015_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_015_src_data),          //          .data
		.out_channel       (width_adapter_015_src_channel),       //          .channel
		.out_valid         (width_adapter_015_src_valid),         //          .valid
		.out_ready         (width_adapter_015_src_ready),         //          .ready
		.out_startofpacket (width_adapter_015_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_016 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src14_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src14_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src14_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src14_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src14_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src14_data),           //          .data
		.out_endofpacket   (width_adapter_016_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_016_src_data),          //          .data
		.out_channel       (width_adapter_016_src_channel),       //          .channel
		.out_valid         (width_adapter_016_src_valid),         //          .valid
		.out_ready         (width_adapter_016_src_ready),         //          .ready
		.out_startofpacket (width_adapter_016_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_017 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_014_src_valid),             //      sink.valid
		.in_channel        (id_router_014_src_channel),           //          .channel
		.in_startofpacket  (id_router_014_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_014_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_014_src_ready),             //          .ready
		.in_data           (id_router_014_src_data),              //          .data
		.out_endofpacket   (width_adapter_017_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_017_src_data),          //          .data
		.out_channel       (width_adapter_017_src_channel),       //          .channel
		.out_valid         (width_adapter_017_src_valid),         //          .valid
		.out_ready         (width_adapter_017_src_ready),         //          .ready
		.out_startofpacket (width_adapter_017_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_018 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src15_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src15_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src15_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src15_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src15_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src15_data),           //          .data
		.out_endofpacket   (width_adapter_018_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_018_src_data),          //          .data
		.out_channel       (width_adapter_018_src_channel),       //          .channel
		.out_valid         (width_adapter_018_src_valid),         //          .valid
		.out_ready         (width_adapter_018_src_ready),         //          .ready
		.out_startofpacket (width_adapter_018_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_019 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_015_src_valid),             //      sink.valid
		.in_channel        (id_router_015_src_channel),           //          .channel
		.in_startofpacket  (id_router_015_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_015_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_015_src_ready),             //          .ready
		.in_data           (id_router_015_src_data),              //          .data
		.out_endofpacket   (width_adapter_019_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_019_src_data),          //          .data
		.out_channel       (width_adapter_019_src_channel),       //          .channel
		.out_valid         (width_adapter_019_src_valid),         //          .valid
		.out_ready         (width_adapter_019_src_ready),         //          .ready
		.out_startofpacket (width_adapter_019_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_020 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src16_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src16_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src16_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src16_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src16_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src16_data),           //          .data
		.out_endofpacket   (width_adapter_020_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_020_src_data),          //          .data
		.out_channel       (width_adapter_020_src_channel),       //          .channel
		.out_valid         (width_adapter_020_src_valid),         //          .valid
		.out_ready         (width_adapter_020_src_ready),         //          .ready
		.out_startofpacket (width_adapter_020_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_021 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_016_src_valid),             //      sink.valid
		.in_channel        (id_router_016_src_channel),           //          .channel
		.in_startofpacket  (id_router_016_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_016_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_016_src_ready),             //          .ready
		.in_data           (id_router_016_src_data),              //          .data
		.out_endofpacket   (width_adapter_021_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_021_src_data),          //          .data
		.out_channel       (width_adapter_021_src_channel),       //          .channel
		.out_valid         (width_adapter_021_src_valid),         //          .valid
		.out_ready         (width_adapter_021_src_ready),         //          .ready
		.out_startofpacket (width_adapter_021_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_022 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src17_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src17_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src17_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src17_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src17_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src17_data),           //          .data
		.out_endofpacket   (width_adapter_022_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_022_src_data),          //          .data
		.out_channel       (width_adapter_022_src_channel),       //          .channel
		.out_valid         (width_adapter_022_src_valid),         //          .valid
		.out_ready         (width_adapter_022_src_ready),         //          .ready
		.out_startofpacket (width_adapter_022_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_023 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_017_src_valid),             //      sink.valid
		.in_channel        (id_router_017_src_channel),           //          .channel
		.in_startofpacket  (id_router_017_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_017_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_017_src_ready),             //          .ready
		.in_data           (id_router_017_src_data),              //          .data
		.out_endofpacket   (width_adapter_023_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_023_src_data),          //          .data
		.out_channel       (width_adapter_023_src_channel),       //          .channel
		.out_valid         (width_adapter_023_src_valid),         //          .valid
		.out_ready         (width_adapter_023_src_ready),         //          .ready
		.out_startofpacket (width_adapter_023_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_024 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src18_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src18_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src18_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src18_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src18_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src18_data),           //          .data
		.out_endofpacket   (width_adapter_024_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_024_src_data),          //          .data
		.out_channel       (width_adapter_024_src_channel),       //          .channel
		.out_valid         (width_adapter_024_src_valid),         //          .valid
		.out_ready         (width_adapter_024_src_ready),         //          .ready
		.out_startofpacket (width_adapter_024_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_025 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_018_src_valid),             //      sink.valid
		.in_channel        (id_router_018_src_channel),           //          .channel
		.in_startofpacket  (id_router_018_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_018_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_018_src_ready),             //          .ready
		.in_data           (id_router_018_src_data),              //          .data
		.out_endofpacket   (width_adapter_025_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_025_src_data),          //          .data
		.out_channel       (width_adapter_025_src_channel),       //          .channel
		.out_valid         (width_adapter_025_src_valid),         //          .valid
		.out_ready         (width_adapter_025_src_ready),         //          .ready
		.out_startofpacket (width_adapter_025_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_026 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src19_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src19_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src19_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src19_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src19_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src19_data),           //          .data
		.out_endofpacket   (width_adapter_026_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_026_src_data),          //          .data
		.out_channel       (width_adapter_026_src_channel),       //          .channel
		.out_valid         (width_adapter_026_src_valid),         //          .valid
		.out_ready         (width_adapter_026_src_ready),         //          .ready
		.out_startofpacket (width_adapter_026_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_027 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_019_src_valid),             //      sink.valid
		.in_channel        (id_router_019_src_channel),           //          .channel
		.in_startofpacket  (id_router_019_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_019_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_019_src_ready),             //          .ready
		.in_data           (id_router_019_src_data),              //          .data
		.out_endofpacket   (width_adapter_027_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_027_src_data),          //          .data
		.out_channel       (width_adapter_027_src_channel),       //          .channel
		.out_valid         (width_adapter_027_src_valid),         //          .valid
		.out_ready         (width_adapter_027_src_ready),         //          .ready
		.out_startofpacket (width_adapter_027_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_028 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src20_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src20_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src20_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src20_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src20_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src20_data),           //          .data
		.out_endofpacket   (width_adapter_028_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_028_src_data),          //          .data
		.out_channel       (width_adapter_028_src_channel),       //          .channel
		.out_valid         (width_adapter_028_src_valid),         //          .valid
		.out_ready         (width_adapter_028_src_ready),         //          .ready
		.out_startofpacket (width_adapter_028_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_029 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_020_src_valid),             //      sink.valid
		.in_channel        (id_router_020_src_channel),           //          .channel
		.in_startofpacket  (id_router_020_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_020_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_020_src_ready),             //          .ready
		.in_data           (id_router_020_src_data),              //          .data
		.out_endofpacket   (width_adapter_029_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_029_src_data),          //          .data
		.out_channel       (width_adapter_029_src_channel),       //          .channel
		.out_valid         (width_adapter_029_src_valid),         //          .valid
		.out_ready         (width_adapter_029_src_ready),         //          .ready
		.out_startofpacket (width_adapter_029_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_030 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src21_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src21_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src21_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src21_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src21_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src21_data),           //          .data
		.out_endofpacket   (width_adapter_030_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_030_src_data),          //          .data
		.out_channel       (width_adapter_030_src_channel),       //          .channel
		.out_valid         (width_adapter_030_src_valid),         //          .valid
		.out_ready         (width_adapter_030_src_ready),         //          .ready
		.out_startofpacket (width_adapter_030_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_031 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_021_src_valid),             //      sink.valid
		.in_channel        (id_router_021_src_channel),           //          .channel
		.in_startofpacket  (id_router_021_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_021_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_021_src_ready),             //          .ready
		.in_data           (id_router_021_src_data),              //          .data
		.out_endofpacket   (width_adapter_031_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_031_src_data),          //          .data
		.out_channel       (width_adapter_031_src_channel),       //          .channel
		.out_valid         (width_adapter_031_src_valid),         //          .valid
		.out_ready         (width_adapter_031_src_ready),         //          .ready
		.out_startofpacket (width_adapter_031_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_032 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src22_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src22_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src22_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src22_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src22_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src22_data),           //          .data
		.out_endofpacket   (width_adapter_032_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_032_src_data),          //          .data
		.out_channel       (width_adapter_032_src_channel),       //          .channel
		.out_valid         (width_adapter_032_src_valid),         //          .valid
		.out_ready         (width_adapter_032_src_ready),         //          .ready
		.out_startofpacket (width_adapter_032_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_033 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_022_src_valid),             //      sink.valid
		.in_channel        (id_router_022_src_channel),           //          .channel
		.in_startofpacket  (id_router_022_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_022_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_022_src_ready),             //          .ready
		.in_data           (id_router_022_src_data),              //          .data
		.out_endofpacket   (width_adapter_033_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_033_src_data),          //          .data
		.out_channel       (width_adapter_033_src_channel),       //          .channel
		.out_valid         (width_adapter_033_src_valid),         //          .valid
		.out_ready         (width_adapter_033_src_ready),         //          .ready
		.out_startofpacket (width_adapter_033_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_034 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src23_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src23_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src23_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src23_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src23_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src23_data),           //          .data
		.out_endofpacket   (width_adapter_034_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_034_src_data),          //          .data
		.out_channel       (width_adapter_034_src_channel),       //          .channel
		.out_valid         (width_adapter_034_src_valid),         //          .valid
		.out_ready         (width_adapter_034_src_ready),         //          .ready
		.out_startofpacket (width_adapter_034_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_035 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_023_src_valid),             //      sink.valid
		.in_channel        (id_router_023_src_channel),           //          .channel
		.in_startofpacket  (id_router_023_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_023_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_023_src_ready),             //          .ready
		.in_data           (id_router_023_src_data),              //          .data
		.out_endofpacket   (width_adapter_035_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_035_src_data),          //          .data
		.out_channel       (width_adapter_035_src_channel),       //          .channel
		.out_valid         (width_adapter_035_src_valid),         //          .valid
		.out_ready         (width_adapter_035_src_ready),         //          .ready
		.out_startofpacket (width_adapter_035_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_036 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src24_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src24_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src24_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src24_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src24_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src24_data),           //          .data
		.out_endofpacket   (width_adapter_036_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_036_src_data),          //          .data
		.out_channel       (width_adapter_036_src_channel),       //          .channel
		.out_valid         (width_adapter_036_src_valid),         //          .valid
		.out_ready         (width_adapter_036_src_ready),         //          .ready
		.out_startofpacket (width_adapter_036_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_037 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_024_src_valid),             //      sink.valid
		.in_channel        (id_router_024_src_channel),           //          .channel
		.in_startofpacket  (id_router_024_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_024_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_024_src_ready),             //          .ready
		.in_data           (id_router_024_src_data),              //          .data
		.out_endofpacket   (width_adapter_037_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_037_src_data),          //          .data
		.out_channel       (width_adapter_037_src_channel),       //          .channel
		.out_valid         (width_adapter_037_src_valid),         //          .valid
		.out_ready         (width_adapter_037_src_ready),         //          .ready
		.out_startofpacket (width_adapter_037_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_038 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src25_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src25_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src25_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src25_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src25_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src25_data),           //          .data
		.out_endofpacket   (width_adapter_038_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_038_src_data),          //          .data
		.out_channel       (width_adapter_038_src_channel),       //          .channel
		.out_valid         (width_adapter_038_src_valid),         //          .valid
		.out_ready         (width_adapter_038_src_ready),         //          .ready
		.out_startofpacket (width_adapter_038_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_039 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_025_src_valid),             //      sink.valid
		.in_channel        (id_router_025_src_channel),           //          .channel
		.in_startofpacket  (id_router_025_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_025_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_025_src_ready),             //          .ready
		.in_data           (id_router_025_src_data),              //          .data
		.out_endofpacket   (width_adapter_039_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_039_src_data),          //          .data
		.out_channel       (width_adapter_039_src_channel),       //          .channel
		.out_valid         (width_adapter_039_src_valid),         //          .valid
		.out_ready         (width_adapter_039_src_ready),         //          .ready
		.out_startofpacket (width_adapter_039_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_040 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src26_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src26_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src26_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src26_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src26_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src26_data),           //          .data
		.out_endofpacket   (width_adapter_040_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_040_src_data),          //          .data
		.out_channel       (width_adapter_040_src_channel),       //          .channel
		.out_valid         (width_adapter_040_src_valid),         //          .valid
		.out_ready         (width_adapter_040_src_ready),         //          .ready
		.out_startofpacket (width_adapter_040_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_041 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_026_src_valid),             //      sink.valid
		.in_channel        (id_router_026_src_channel),           //          .channel
		.in_startofpacket  (id_router_026_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_026_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_026_src_ready),             //          .ready
		.in_data           (id_router_026_src_data),              //          .data
		.out_endofpacket   (width_adapter_041_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_041_src_data),          //          .data
		.out_channel       (width_adapter_041_src_channel),       //          .channel
		.out_valid         (width_adapter_041_src_valid),         //          .valid
		.out_ready         (width_adapter_041_src_ready),         //          .ready
		.out_startofpacket (width_adapter_041_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_042 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src27_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src27_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src27_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src27_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src27_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src27_data),           //          .data
		.out_endofpacket   (width_adapter_042_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_042_src_data),          //          .data
		.out_channel       (width_adapter_042_src_channel),       //          .channel
		.out_valid         (width_adapter_042_src_valid),         //          .valid
		.out_ready         (width_adapter_042_src_ready),         //          .ready
		.out_startofpacket (width_adapter_042_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_043 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_027_src_valid),             //      sink.valid
		.in_channel        (id_router_027_src_channel),           //          .channel
		.in_startofpacket  (id_router_027_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_027_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_027_src_ready),             //          .ready
		.in_data           (id_router_027_src_data),              //          .data
		.out_endofpacket   (width_adapter_043_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_043_src_data),          //          .data
		.out_channel       (width_adapter_043_src_channel),       //          .channel
		.out_valid         (width_adapter_043_src_valid),         //          .valid
		.out_ready         (width_adapter_043_src_ready),         //          .ready
		.out_startofpacket (width_adapter_043_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_044 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src28_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src28_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src28_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src28_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src28_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src28_data),           //          .data
		.out_endofpacket   (width_adapter_044_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_044_src_data),          //          .data
		.out_channel       (width_adapter_044_src_channel),       //          .channel
		.out_valid         (width_adapter_044_src_valid),         //          .valid
		.out_ready         (width_adapter_044_src_ready),         //          .ready
		.out_startofpacket (width_adapter_044_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_045 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_028_src_valid),             //      sink.valid
		.in_channel        (id_router_028_src_channel),           //          .channel
		.in_startofpacket  (id_router_028_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_028_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_028_src_ready),             //          .ready
		.in_data           (id_router_028_src_data),              //          .data
		.out_endofpacket   (width_adapter_045_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_045_src_data),          //          .data
		.out_channel       (width_adapter_045_src_channel),       //          .channel
		.out_valid         (width_adapter_045_src_valid),         //          .valid
		.out_ready         (width_adapter_045_src_ready),         //          .ready
		.out_startofpacket (width_adapter_045_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_046 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src29_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src29_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src29_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src29_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src29_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src29_data),           //          .data
		.out_endofpacket   (width_adapter_046_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_046_src_data),          //          .data
		.out_channel       (width_adapter_046_src_channel),       //          .channel
		.out_valid         (width_adapter_046_src_valid),         //          .valid
		.out_ready         (width_adapter_046_src_ready),         //          .ready
		.out_startofpacket (width_adapter_046_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_047 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_029_src_valid),             //      sink.valid
		.in_channel        (id_router_029_src_channel),           //          .channel
		.in_startofpacket  (id_router_029_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_029_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_029_src_ready),             //          .ready
		.in_data           (id_router_029_src_data),              //          .data
		.out_endofpacket   (width_adapter_047_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_047_src_data),          //          .data
		.out_channel       (width_adapter_047_src_channel),       //          .channel
		.out_valid         (width_adapter_047_src_valid),         //          .valid
		.out_ready         (width_adapter_047_src_ready),         //          .ready
		.out_startofpacket (width_adapter_047_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_048 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src30_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src30_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src30_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src30_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src30_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src30_data),           //          .data
		.out_endofpacket   (width_adapter_048_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_048_src_data),          //          .data
		.out_channel       (width_adapter_048_src_channel),       //          .channel
		.out_valid         (width_adapter_048_src_valid),         //          .valid
		.out_ready         (width_adapter_048_src_ready),         //          .ready
		.out_startofpacket (width_adapter_048_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_049 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_030_src_valid),             //      sink.valid
		.in_channel        (id_router_030_src_channel),           //          .channel
		.in_startofpacket  (id_router_030_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_030_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_030_src_ready),             //          .ready
		.in_data           (id_router_030_src_data),              //          .data
		.out_endofpacket   (width_adapter_049_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_049_src_data),          //          .data
		.out_channel       (width_adapter_049_src_channel),       //          .channel
		.out_valid         (width_adapter_049_src_valid),         //          .valid
		.out_ready         (width_adapter_049_src_ready),         //          .ready
		.out_startofpacket (width_adapter_049_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_050 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src31_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src31_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src31_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src31_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src31_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src31_data),           //          .data
		.out_endofpacket   (width_adapter_050_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_050_src_data),          //          .data
		.out_channel       (width_adapter_050_src_channel),       //          .channel
		.out_valid         (width_adapter_050_src_valid),         //          .valid
		.out_ready         (width_adapter_050_src_ready),         //          .ready
		.out_startofpacket (width_adapter_050_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_051 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_031_src_valid),             //      sink.valid
		.in_channel        (id_router_031_src_channel),           //          .channel
		.in_startofpacket  (id_router_031_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_031_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_031_src_ready),             //          .ready
		.in_data           (id_router_031_src_data),              //          .data
		.out_endofpacket   (width_adapter_051_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_051_src_data),          //          .data
		.out_channel       (width_adapter_051_src_channel),       //          .channel
		.out_valid         (width_adapter_051_src_valid),         //          .valid
		.out_ready         (width_adapter_051_src_ready),         //          .ready
		.out_startofpacket (width_adapter_051_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_052 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src32_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src32_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src32_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src32_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src32_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src32_data),           //          .data
		.out_endofpacket   (width_adapter_052_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_052_src_data),          //          .data
		.out_channel       (width_adapter_052_src_channel),       //          .channel
		.out_valid         (width_adapter_052_src_valid),         //          .valid
		.out_ready         (width_adapter_052_src_ready),         //          .ready
		.out_startofpacket (width_adapter_052_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_053 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_032_src_valid),             //      sink.valid
		.in_channel        (id_router_032_src_channel),           //          .channel
		.in_startofpacket  (id_router_032_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_032_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_032_src_ready),             //          .ready
		.in_data           (id_router_032_src_data),              //          .data
		.out_endofpacket   (width_adapter_053_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_053_src_data),          //          .data
		.out_channel       (width_adapter_053_src_channel),       //          .channel
		.out_valid         (width_adapter_053_src_valid),         //          .valid
		.out_ready         (width_adapter_053_src_ready),         //          .ready
		.out_startofpacket (width_adapter_053_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_054 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src33_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src33_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src33_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src33_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src33_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src33_data),           //          .data
		.out_endofpacket   (width_adapter_054_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_054_src_data),          //          .data
		.out_channel       (width_adapter_054_src_channel),       //          .channel
		.out_valid         (width_adapter_054_src_valid),         //          .valid
		.out_ready         (width_adapter_054_src_ready),         //          .ready
		.out_startofpacket (width_adapter_054_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_055 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_033_src_valid),             //      sink.valid
		.in_channel        (id_router_033_src_channel),           //          .channel
		.in_startofpacket  (id_router_033_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_033_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_033_src_ready),             //          .ready
		.in_data           (id_router_033_src_data),              //          .data
		.out_endofpacket   (width_adapter_055_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_055_src_data),          //          .data
		.out_channel       (width_adapter_055_src_channel),       //          .channel
		.out_valid         (width_adapter_055_src_valid),         //          .valid
		.out_ready         (width_adapter_055_src_ready),         //          .ready
		.out_startofpacket (width_adapter_055_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_056 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src34_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src34_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src34_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src34_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src34_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src34_data),           //          .data
		.out_endofpacket   (width_adapter_056_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_056_src_data),          //          .data
		.out_channel       (width_adapter_056_src_channel),       //          .channel
		.out_valid         (width_adapter_056_src_valid),         //          .valid
		.out_ready         (width_adapter_056_src_ready),         //          .ready
		.out_startofpacket (width_adapter_056_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_057 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_034_src_valid),             //      sink.valid
		.in_channel        (id_router_034_src_channel),           //          .channel
		.in_startofpacket  (id_router_034_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_034_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_034_src_ready),             //          .ready
		.in_data           (id_router_034_src_data),              //          .data
		.out_endofpacket   (width_adapter_057_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_057_src_data),          //          .data
		.out_channel       (width_adapter_057_src_channel),       //          .channel
		.out_valid         (width_adapter_057_src_valid),         //          .valid
		.out_ready         (width_adapter_057_src_ready),         //          .ready
		.out_startofpacket (width_adapter_057_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_058 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src35_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src35_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src35_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src35_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src35_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src35_data),           //          .data
		.out_endofpacket   (width_adapter_058_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_058_src_data),          //          .data
		.out_channel       (width_adapter_058_src_channel),       //          .channel
		.out_valid         (width_adapter_058_src_valid),         //          .valid
		.out_ready         (width_adapter_058_src_ready),         //          .ready
		.out_startofpacket (width_adapter_058_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_059 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_035_src_valid),             //      sink.valid
		.in_channel        (id_router_035_src_channel),           //          .channel
		.in_startofpacket  (id_router_035_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_035_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_035_src_ready),             //          .ready
		.in_data           (id_router_035_src_data),              //          .data
		.out_endofpacket   (width_adapter_059_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_059_src_data),          //          .data
		.out_channel       (width_adapter_059_src_channel),       //          .channel
		.out_valid         (width_adapter_059_src_valid),         //          .valid
		.out_ready         (width_adapter_059_src_ready),         //          .ready
		.out_startofpacket (width_adapter_059_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_060 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src36_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src36_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src36_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src36_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src36_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src36_data),           //          .data
		.out_endofpacket   (width_adapter_060_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_060_src_data),          //          .data
		.out_channel       (width_adapter_060_src_channel),       //          .channel
		.out_valid         (width_adapter_060_src_valid),         //          .valid
		.out_ready         (width_adapter_060_src_ready),         //          .ready
		.out_startofpacket (width_adapter_060_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_061 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_036_src_valid),             //      sink.valid
		.in_channel        (id_router_036_src_channel),           //          .channel
		.in_startofpacket  (id_router_036_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_036_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_036_src_ready),             //          .ready
		.in_data           (id_router_036_src_data),              //          .data
		.out_endofpacket   (width_adapter_061_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_061_src_data),          //          .data
		.out_channel       (width_adapter_061_src_channel),       //          .channel
		.out_valid         (width_adapter_061_src_valid),         //          .valid
		.out_ready         (width_adapter_061_src_ready),         //          .ready
		.out_startofpacket (width_adapter_061_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_062 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src37_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src37_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src37_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src37_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src37_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src37_data),           //          .data
		.out_endofpacket   (width_adapter_062_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_062_src_data),          //          .data
		.out_channel       (width_adapter_062_src_channel),       //          .channel
		.out_valid         (width_adapter_062_src_valid),         //          .valid
		.out_ready         (width_adapter_062_src_ready),         //          .ready
		.out_startofpacket (width_adapter_062_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_063 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_037_src_valid),             //      sink.valid
		.in_channel        (id_router_037_src_channel),           //          .channel
		.in_startofpacket  (id_router_037_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_037_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_037_src_ready),             //          .ready
		.in_data           (id_router_037_src_data),              //          .data
		.out_endofpacket   (width_adapter_063_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_063_src_data),          //          .data
		.out_channel       (width_adapter_063_src_channel),       //          .channel
		.out_valid         (width_adapter_063_src_valid),         //          .valid
		.out_ready         (width_adapter_063_src_ready),         //          .ready
		.out_startofpacket (width_adapter_063_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_064 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src38_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src38_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src38_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src38_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src38_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src38_data),           //          .data
		.out_endofpacket   (width_adapter_064_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_064_src_data),          //          .data
		.out_channel       (width_adapter_064_src_channel),       //          .channel
		.out_valid         (width_adapter_064_src_valid),         //          .valid
		.out_ready         (width_adapter_064_src_ready),         //          .ready
		.out_startofpacket (width_adapter_064_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_065 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_038_src_valid),             //      sink.valid
		.in_channel        (id_router_038_src_channel),           //          .channel
		.in_startofpacket  (id_router_038_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_038_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_038_src_ready),             //          .ready
		.in_data           (id_router_038_src_data),              //          .data
		.out_endofpacket   (width_adapter_065_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_065_src_data),          //          .data
		.out_channel       (width_adapter_065_src_channel),       //          .channel
		.out_valid         (width_adapter_065_src_valid),         //          .valid
		.out_ready         (width_adapter_065_src_ready),         //          .ready
		.out_startofpacket (width_adapter_065_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_066 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src39_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src39_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src39_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src39_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src39_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src39_data),           //          .data
		.out_endofpacket   (width_adapter_066_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_066_src_data),          //          .data
		.out_channel       (width_adapter_066_src_channel),       //          .channel
		.out_valid         (width_adapter_066_src_valid),         //          .valid
		.out_ready         (width_adapter_066_src_ready),         //          .ready
		.out_startofpacket (width_adapter_066_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_067 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_039_src_valid),             //      sink.valid
		.in_channel        (id_router_039_src_channel),           //          .channel
		.in_startofpacket  (id_router_039_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_039_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_039_src_ready),             //          .ready
		.in_data           (id_router_039_src_data),              //          .data
		.out_endofpacket   (width_adapter_067_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_067_src_data),          //          .data
		.out_channel       (width_adapter_067_src_channel),       //          .channel
		.out_valid         (width_adapter_067_src_valid),         //          .valid
		.out_ready         (width_adapter_067_src_ready),         //          .ready
		.out_startofpacket (width_adapter_067_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_068 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src40_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src40_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src40_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src40_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src40_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src40_data),           //          .data
		.out_endofpacket   (width_adapter_068_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_068_src_data),          //          .data
		.out_channel       (width_adapter_068_src_channel),       //          .channel
		.out_valid         (width_adapter_068_src_valid),         //          .valid
		.out_ready         (width_adapter_068_src_ready),         //          .ready
		.out_startofpacket (width_adapter_068_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_069 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_040_src_valid),             //      sink.valid
		.in_channel        (id_router_040_src_channel),           //          .channel
		.in_startofpacket  (id_router_040_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_040_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_040_src_ready),             //          .ready
		.in_data           (id_router_040_src_data),              //          .data
		.out_endofpacket   (width_adapter_069_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_069_src_data),          //          .data
		.out_channel       (width_adapter_069_src_channel),       //          .channel
		.out_valid         (width_adapter_069_src_valid),         //          .valid
		.out_ready         (width_adapter_069_src_ready),         //          .ready
		.out_startofpacket (width_adapter_069_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_070 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src41_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src41_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src41_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src41_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src41_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src41_data),           //          .data
		.out_endofpacket   (width_adapter_070_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_070_src_data),          //          .data
		.out_channel       (width_adapter_070_src_channel),       //          .channel
		.out_valid         (width_adapter_070_src_valid),         //          .valid
		.out_ready         (width_adapter_070_src_ready),         //          .ready
		.out_startofpacket (width_adapter_070_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_071 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_041_src_valid),             //      sink.valid
		.in_channel        (id_router_041_src_channel),           //          .channel
		.in_startofpacket  (id_router_041_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_041_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_041_src_ready),             //          .ready
		.in_data           (id_router_041_src_data),              //          .data
		.out_endofpacket   (width_adapter_071_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_071_src_data),          //          .data
		.out_channel       (width_adapter_071_src_channel),       //          .channel
		.out_valid         (width_adapter_071_src_valid),         //          .valid
		.out_ready         (width_adapter_071_src_ready),         //          .ready
		.out_startofpacket (width_adapter_071_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_072 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src42_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src42_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src42_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src42_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src42_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src42_data),           //          .data
		.out_endofpacket   (width_adapter_072_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_072_src_data),          //          .data
		.out_channel       (width_adapter_072_src_channel),       //          .channel
		.out_valid         (width_adapter_072_src_valid),         //          .valid
		.out_ready         (width_adapter_072_src_ready),         //          .ready
		.out_startofpacket (width_adapter_072_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_073 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_042_src_valid),             //      sink.valid
		.in_channel        (id_router_042_src_channel),           //          .channel
		.in_startofpacket  (id_router_042_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_042_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_042_src_ready),             //          .ready
		.in_data           (id_router_042_src_data),              //          .data
		.out_endofpacket   (width_adapter_073_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_073_src_data),          //          .data
		.out_channel       (width_adapter_073_src_channel),       //          .channel
		.out_valid         (width_adapter_073_src_valid),         //          .valid
		.out_ready         (width_adapter_073_src_ready),         //          .ready
		.out_startofpacket (width_adapter_073_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_074 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src43_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src43_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src43_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src43_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src43_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src43_data),           //          .data
		.out_endofpacket   (width_adapter_074_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_074_src_data),          //          .data
		.out_channel       (width_adapter_074_src_channel),       //          .channel
		.out_valid         (width_adapter_074_src_valid),         //          .valid
		.out_ready         (width_adapter_074_src_ready),         //          .ready
		.out_startofpacket (width_adapter_074_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_075 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_043_src_valid),             //      sink.valid
		.in_channel        (id_router_043_src_channel),           //          .channel
		.in_startofpacket  (id_router_043_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_043_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_043_src_ready),             //          .ready
		.in_data           (id_router_043_src_data),              //          .data
		.out_endofpacket   (width_adapter_075_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_075_src_data),          //          .data
		.out_channel       (width_adapter_075_src_channel),       //          .channel
		.out_valid         (width_adapter_075_src_valid),         //          .valid
		.out_ready         (width_adapter_075_src_ready),         //          .ready
		.out_startofpacket (width_adapter_075_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_076 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src44_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src44_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src44_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src44_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src44_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src44_data),           //          .data
		.out_endofpacket   (width_adapter_076_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_076_src_data),          //          .data
		.out_channel       (width_adapter_076_src_channel),       //          .channel
		.out_valid         (width_adapter_076_src_valid),         //          .valid
		.out_ready         (width_adapter_076_src_ready),         //          .ready
		.out_startofpacket (width_adapter_076_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_077 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_044_src_valid),             //      sink.valid
		.in_channel        (id_router_044_src_channel),           //          .channel
		.in_startofpacket  (id_router_044_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_044_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_044_src_ready),             //          .ready
		.in_data           (id_router_044_src_data),              //          .data
		.out_endofpacket   (width_adapter_077_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_077_src_data),          //          .data
		.out_channel       (width_adapter_077_src_channel),       //          .channel
		.out_valid         (width_adapter_077_src_valid),         //          .valid
		.out_ready         (width_adapter_077_src_ready),         //          .ready
		.out_startofpacket (width_adapter_077_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_078 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src45_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src45_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src45_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src45_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src45_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src45_data),           //          .data
		.out_endofpacket   (width_adapter_078_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_078_src_data),          //          .data
		.out_channel       (width_adapter_078_src_channel),       //          .channel
		.out_valid         (width_adapter_078_src_valid),         //          .valid
		.out_ready         (width_adapter_078_src_ready),         //          .ready
		.out_startofpacket (width_adapter_078_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_079 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_045_src_valid),             //      sink.valid
		.in_channel        (id_router_045_src_channel),           //          .channel
		.in_startofpacket  (id_router_045_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_045_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_045_src_ready),             //          .ready
		.in_data           (id_router_045_src_data),              //          .data
		.out_endofpacket   (width_adapter_079_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_079_src_data),          //          .data
		.out_channel       (width_adapter_079_src_channel),       //          .channel
		.out_valid         (width_adapter_079_src_valid),         //          .valid
		.out_ready         (width_adapter_079_src_ready),         //          .ready
		.out_startofpacket (width_adapter_079_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_080 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src46_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src46_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src46_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src46_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src46_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src46_data),           //          .data
		.out_endofpacket   (width_adapter_080_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_080_src_data),          //          .data
		.out_channel       (width_adapter_080_src_channel),       //          .channel
		.out_valid         (width_adapter_080_src_valid),         //          .valid
		.out_ready         (width_adapter_080_src_ready),         //          .ready
		.out_startofpacket (width_adapter_080_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_081 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_046_src_valid),             //      sink.valid
		.in_channel        (id_router_046_src_channel),           //          .channel
		.in_startofpacket  (id_router_046_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_046_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_046_src_ready),             //          .ready
		.in_data           (id_router_046_src_data),              //          .data
		.out_endofpacket   (width_adapter_081_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_081_src_data),          //          .data
		.out_channel       (width_adapter_081_src_channel),       //          .channel
		.out_valid         (width_adapter_081_src_valid),         //          .valid
		.out_ready         (width_adapter_081_src_ready),         //          .ready
		.out_startofpacket (width_adapter_081_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_082 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src47_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src47_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src47_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src47_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src47_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src47_data),           //          .data
		.out_endofpacket   (width_adapter_082_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_082_src_data),          //          .data
		.out_channel       (width_adapter_082_src_channel),       //          .channel
		.out_valid         (width_adapter_082_src_valid),         //          .valid
		.out_ready         (width_adapter_082_src_ready),         //          .ready
		.out_startofpacket (width_adapter_082_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_083 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_047_src_valid),             //      sink.valid
		.in_channel        (id_router_047_src_channel),           //          .channel
		.in_startofpacket  (id_router_047_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_047_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_047_src_ready),             //          .ready
		.in_data           (id_router_047_src_data),              //          .data
		.out_endofpacket   (width_adapter_083_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_083_src_data),          //          .data
		.out_channel       (width_adapter_083_src_channel),       //          .channel
		.out_valid         (width_adapter_083_src_valid),         //          .valid
		.out_ready         (width_adapter_083_src_ready),         //          .ready
		.out_startofpacket (width_adapter_083_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_084 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src48_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src48_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src48_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src48_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src48_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src48_data),           //          .data
		.out_endofpacket   (width_adapter_084_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_084_src_data),          //          .data
		.out_channel       (width_adapter_084_src_channel),       //          .channel
		.out_valid         (width_adapter_084_src_valid),         //          .valid
		.out_ready         (width_adapter_084_src_ready),         //          .ready
		.out_startofpacket (width_adapter_084_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_085 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_048_src_valid),             //      sink.valid
		.in_channel        (id_router_048_src_channel),           //          .channel
		.in_startofpacket  (id_router_048_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_048_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_048_src_ready),             //          .ready
		.in_data           (id_router_048_src_data),              //          .data
		.out_endofpacket   (width_adapter_085_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_085_src_data),          //          .data
		.out_channel       (width_adapter_085_src_channel),       //          .channel
		.out_valid         (width_adapter_085_src_valid),         //          .valid
		.out_ready         (width_adapter_085_src_ready),         //          .ready
		.out_startofpacket (width_adapter_085_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_086 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src49_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src49_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src49_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src49_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src49_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src49_data),           //          .data
		.out_endofpacket   (width_adapter_086_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_086_src_data),          //          .data
		.out_channel       (width_adapter_086_src_channel),       //          .channel
		.out_valid         (width_adapter_086_src_valid),         //          .valid
		.out_ready         (width_adapter_086_src_ready),         //          .ready
		.out_startofpacket (width_adapter_086_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_087 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_049_src_valid),             //      sink.valid
		.in_channel        (id_router_049_src_channel),           //          .channel
		.in_startofpacket  (id_router_049_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_049_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_049_src_ready),             //          .ready
		.in_data           (id_router_049_src_data),              //          .data
		.out_endofpacket   (width_adapter_087_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_087_src_data),          //          .data
		.out_channel       (width_adapter_087_src_channel),       //          .channel
		.out_valid         (width_adapter_087_src_valid),         //          .valid
		.out_ready         (width_adapter_087_src_ready),         //          .ready
		.out_startofpacket (width_adapter_087_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_088 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src50_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src50_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src50_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src50_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src50_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src50_data),           //          .data
		.out_endofpacket   (width_adapter_088_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_088_src_data),          //          .data
		.out_channel       (width_adapter_088_src_channel),       //          .channel
		.out_valid         (width_adapter_088_src_valid),         //          .valid
		.out_ready         (width_adapter_088_src_ready),         //          .ready
		.out_startofpacket (width_adapter_088_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_089 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_050_src_valid),             //      sink.valid
		.in_channel        (id_router_050_src_channel),           //          .channel
		.in_startofpacket  (id_router_050_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_050_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_050_src_ready),             //          .ready
		.in_data           (id_router_050_src_data),              //          .data
		.out_endofpacket   (width_adapter_089_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_089_src_data),          //          .data
		.out_channel       (width_adapter_089_src_channel),       //          .channel
		.out_valid         (width_adapter_089_src_valid),         //          .valid
		.out_ready         (width_adapter_089_src_ready),         //          .ready
		.out_startofpacket (width_adapter_089_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_090 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src51_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src51_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src51_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src51_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src51_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src51_data),           //          .data
		.out_endofpacket   (width_adapter_090_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_090_src_data),          //          .data
		.out_channel       (width_adapter_090_src_channel),       //          .channel
		.out_valid         (width_adapter_090_src_valid),         //          .valid
		.out_ready         (width_adapter_090_src_ready),         //          .ready
		.out_startofpacket (width_adapter_090_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_091 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_051_src_valid),             //      sink.valid
		.in_channel        (id_router_051_src_channel),           //          .channel
		.in_startofpacket  (id_router_051_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_051_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_051_src_ready),             //          .ready
		.in_data           (id_router_051_src_data),              //          .data
		.out_endofpacket   (width_adapter_091_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_091_src_data),          //          .data
		.out_channel       (width_adapter_091_src_channel),       //          .channel
		.out_valid         (width_adapter_091_src_valid),         //          .valid
		.out_ready         (width_adapter_091_src_ready),         //          .ready
		.out_startofpacket (width_adapter_091_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_092 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src52_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src52_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src52_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src52_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src52_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src52_data),           //          .data
		.out_endofpacket   (width_adapter_092_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_092_src_data),          //          .data
		.out_channel       (width_adapter_092_src_channel),       //          .channel
		.out_valid         (width_adapter_092_src_valid),         //          .valid
		.out_ready         (width_adapter_092_src_ready),         //          .ready
		.out_startofpacket (width_adapter_092_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_093 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_052_src_valid),             //      sink.valid
		.in_channel        (id_router_052_src_channel),           //          .channel
		.in_startofpacket  (id_router_052_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_052_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_052_src_ready),             //          .ready
		.in_data           (id_router_052_src_data),              //          .data
		.out_endofpacket   (width_adapter_093_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_093_src_data),          //          .data
		.out_channel       (width_adapter_093_src_channel),       //          .channel
		.out_valid         (width_adapter_093_src_valid),         //          .valid
		.out_ready         (width_adapter_093_src_ready),         //          .ready
		.out_startofpacket (width_adapter_093_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_094 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src53_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src53_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src53_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src53_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src53_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src53_data),           //          .data
		.out_endofpacket   (width_adapter_094_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_094_src_data),          //          .data
		.out_channel       (width_adapter_094_src_channel),       //          .channel
		.out_valid         (width_adapter_094_src_valid),         //          .valid
		.out_ready         (width_adapter_094_src_ready),         //          .ready
		.out_startofpacket (width_adapter_094_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_095 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_053_src_valid),             //      sink.valid
		.in_channel        (id_router_053_src_channel),           //          .channel
		.in_startofpacket  (id_router_053_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_053_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_053_src_ready),             //          .ready
		.in_data           (id_router_053_src_data),              //          .data
		.out_endofpacket   (width_adapter_095_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_095_src_data),          //          .data
		.out_channel       (width_adapter_095_src_channel),       //          .channel
		.out_valid         (width_adapter_095_src_valid),         //          .valid
		.out_ready         (width_adapter_095_src_ready),         //          .ready
		.out_startofpacket (width_adapter_095_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_096 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src54_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src54_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src54_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src54_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src54_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src54_data),           //          .data
		.out_endofpacket   (width_adapter_096_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_096_src_data),          //          .data
		.out_channel       (width_adapter_096_src_channel),       //          .channel
		.out_valid         (width_adapter_096_src_valid),         //          .valid
		.out_ready         (width_adapter_096_src_ready),         //          .ready
		.out_startofpacket (width_adapter_096_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_097 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_054_src_valid),             //      sink.valid
		.in_channel        (id_router_054_src_channel),           //          .channel
		.in_startofpacket  (id_router_054_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_054_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_054_src_ready),             //          .ready
		.in_data           (id_router_054_src_data),              //          .data
		.out_endofpacket   (width_adapter_097_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_097_src_data),          //          .data
		.out_channel       (width_adapter_097_src_channel),       //          .channel
		.out_valid         (width_adapter_097_src_valid),         //          .valid
		.out_ready         (width_adapter_097_src_ready),         //          .ready
		.out_startofpacket (width_adapter_097_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_098 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src55_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src55_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src55_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src55_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src55_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src55_data),           //          .data
		.out_endofpacket   (width_adapter_098_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_098_src_data),          //          .data
		.out_channel       (width_adapter_098_src_channel),       //          .channel
		.out_valid         (width_adapter_098_src_valid),         //          .valid
		.out_ready         (width_adapter_098_src_ready),         //          .ready
		.out_startofpacket (width_adapter_098_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_099 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_055_src_valid),             //      sink.valid
		.in_channel        (id_router_055_src_channel),           //          .channel
		.in_startofpacket  (id_router_055_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_055_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_055_src_ready),             //          .ready
		.in_data           (id_router_055_src_data),              //          .data
		.out_endofpacket   (width_adapter_099_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_099_src_data),          //          .data
		.out_channel       (width_adapter_099_src_channel),       //          .channel
		.out_valid         (width_adapter_099_src_valid),         //          .valid
		.out_ready         (width_adapter_099_src_ready),         //          .ready
		.out_startofpacket (width_adapter_099_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_100 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src56_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src56_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src56_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src56_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src56_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src56_data),           //          .data
		.out_endofpacket   (width_adapter_100_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_100_src_data),          //          .data
		.out_channel       (width_adapter_100_src_channel),       //          .channel
		.out_valid         (width_adapter_100_src_valid),         //          .valid
		.out_ready         (width_adapter_100_src_ready),         //          .ready
		.out_startofpacket (width_adapter_100_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_101 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_056_src_valid),             //      sink.valid
		.in_channel        (id_router_056_src_channel),           //          .channel
		.in_startofpacket  (id_router_056_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_056_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_056_src_ready),             //          .ready
		.in_data           (id_router_056_src_data),              //          .data
		.out_endofpacket   (width_adapter_101_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_101_src_data),          //          .data
		.out_channel       (width_adapter_101_src_channel),       //          .channel
		.out_valid         (width_adapter_101_src_valid),         //          .valid
		.out_ready         (width_adapter_101_src_ready),         //          .ready
		.out_startofpacket (width_adapter_101_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (75),
		.IN_PKT_BYTE_CNT_L             (73),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (78),
		.IN_PKT_BURSTWRAP_L            (76),
		.IN_ST_DATA_W                  (93),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (48),
		.OUT_PKT_BYTE_CNT_L            (46),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_ST_DATA_W                 (66),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_102 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (cmd_xbar_demux_src57_valid),          //      sink.valid
		.in_channel        (cmd_xbar_demux_src57_channel),        //          .channel
		.in_startofpacket  (cmd_xbar_demux_src57_startofpacket),  //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src57_endofpacket),    //          .endofpacket
		.in_ready          (cmd_xbar_demux_src57_ready),          //          .ready
		.in_data           (cmd_xbar_demux_src57_data),           //          .data
		.out_endofpacket   (width_adapter_102_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_102_src_data),          //          .data
		.out_channel       (width_adapter_102_src_channel),       //          .channel
		.out_valid         (width_adapter_102_src_valid),         //          .valid
		.out_ready         (width_adapter_102_src_ready),         //          .ready
		.out_startofpacket (width_adapter_102_src_startofpacket)  //          .startofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (48),
		.IN_PKT_BYTE_CNT_L             (46),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (51),
		.IN_PKT_BURSTWRAP_L            (49),
		.IN_ST_DATA_W                  (66),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (75),
		.OUT_PKT_BYTE_CNT_L            (73),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_ST_DATA_W                 (93),
		.ST_CHANNEL_W                  (58),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_103 (
		.clk               (sam9_mclk_clk),                       //       clk.clk
		.reset             (sam9_mrst_reset),                     // clk_reset.reset
		.in_valid          (id_router_057_src_valid),             //      sink.valid
		.in_channel        (id_router_057_src_channel),           //          .channel
		.in_startofpacket  (id_router_057_src_startofpacket),     //          .startofpacket
		.in_endofpacket    (id_router_057_src_endofpacket),       //          .endofpacket
		.in_ready          (id_router_057_src_ready),             //          .ready
		.in_data           (id_router_057_src_data),              //          .data
		.out_endofpacket   (width_adapter_103_src_endofpacket),   //       src.endofpacket
		.out_data          (width_adapter_103_src_data),          //          .data
		.out_channel       (width_adapter_103_src_channel),       //          .channel
		.out_valid         (width_adapter_103_src_valid),         //          .valid
		.out_ready         (width_adapter_103_src_ready),         //          .ready
		.out_startofpacket (width_adapter_103_src_startofpacket)  //          .startofpacket
	);

	frontier_irq_mapper irq_mapper (
		.clk           (sam9_mclk_clk),                 //       clk.clk
		.reset         (sam9_mrst_reset),               // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),      // receiver0.irq
		.sender_irq    (irq_synchronizer_receiver_irq)  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (10)
	) irq_synchronizer (
		.receiver_clk   (sam9_mclk_clk),                 //       receiver_clk.clk
		.sender_clk     (sam9_mclk_clk),                 //         sender_clk.clk
		.receiver_reset (sam9_mrst_reset),               // receiver_clk_reset.reset
		.sender_reset   (sam9_mrst_reset),               //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq), //           receiver.irq
		.sender_irq     (sam9_events_irq)                //             sender.irq
	);

endmodule
