// frontier.v

// Generated using ACDS version 11.1sp2 259 at 2012.07.22.11:10:12

`timescale 1 ps / 1 ps
module frontier (
		input  wire        m1_RSTN,  // m1.RSTN
		input  wire        m1_CLK,   //   .CLK
		input  wire [21:0] m1_ADDR,  //   .ADDR
		inout  wire [31:0] m1_DATA,  //   .DATA
		input  wire [3:0]  m1_CSN,   //   .CSN
		input  wire [3:0]  m1_BEN,   //   .BEN
		input  wire        m1_RDN,   //   .RDN
		input  wire        m1_WRN,   //   .WRN
		output wire        m1_WAITN, //   .WAITN
		output wire [9:0]  m1_EINT   //   .EINT
	);

	wire         hps_tabby_mrst_reset;                                                                         // HPS_Tabby:rso_MRST_reset -> [HPS_Tabby_M1_translator:reset, HPS_Tabby_M1_translator_avalon_universal_master_0_agent:reset, SysID:rsi_MRST_reset, SysID_SysID_translator:reset, SysID_SysID_translator_avalon_universal_slave_0_agent:reset, SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, cmd_xbar_demux:reset, id_router:reset, id_router_001:reset, irq_mapper:reset, irq_synchronizer:receiver_reset, irq_synchronizer:sender_reset, limiter:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_mux:reset, test_RegWaitRW32_0:rsi_MRST_reset, test_RegWaitRW32_0_test_translator:reset, test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:reset, test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         hps_tabby_mclk_clk;                                                                           // HPS_Tabby:cso_MCLK_clk -> [HPS_Tabby_M1_translator:clk, HPS_Tabby_M1_translator_avalon_universal_master_0_agent:clk, SysID:csi_MCLK_clk, SysID_SysID_translator:clk, SysID_SysID_translator_avalon_universal_slave_0_agent:clk, SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, cmd_xbar_demux:clk, id_router:clk, id_router_001:clk, irq_mapper:clk, irq_synchronizer:receiver_clk, irq_synchronizer:sender_clk, limiter:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_mux:clk, test_RegWaitRW32_0:csi_MCLK_clk, test_RegWaitRW32_0_test_translator:clk, test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:clk, test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire         hps_tabby_m1_waitrequest;                                                                     // HPS_Tabby_M1_translator:av_waitrequest -> HPS_Tabby:avm_M1_waitrequest
	wire  [29:0] hps_tabby_m1_address;                                                                         // HPS_Tabby:avm_M1_address -> HPS_Tabby_M1_translator:av_address
	wire  [31:0] hps_tabby_m1_writedata;                                                                       // HPS_Tabby:avm_M1_writedata -> HPS_Tabby_M1_translator:av_writedata
	wire         hps_tabby_m1_write;                                                                           // HPS_Tabby:avm_M1_write -> HPS_Tabby_M1_translator:av_write
	wire         hps_tabby_m1_read;                                                                            // HPS_Tabby:avm_M1_read -> HPS_Tabby_M1_translator:av_read
	wire  [31:0] hps_tabby_m1_readdata;                                                                        // HPS_Tabby_M1_translator:av_readdata -> HPS_Tabby:avm_M1_readdata
	wire         hps_tabby_m1_begintransfer;                                                                   // HPS_Tabby:avm_M1_begintransfer -> HPS_Tabby_M1_translator:av_begintransfer
	wire         hps_tabby_m1_readdatavalid;                                                                   // HPS_Tabby_M1_translator:av_readdatavalid -> HPS_Tabby:avm_M1_readdatavalid
	wire   [3:0] hps_tabby_m1_byteenable;                                                                      // HPS_Tabby:avm_M1_byteenable -> HPS_Tabby_M1_translator:av_byteenable
	wire         sysid_sysid_translator_avalon_anti_slave_0_waitrequest;                                       // SysID:avs_SysID_waitrequest -> SysID_SysID_translator:av_waitrequest
	wire   [1:0] sysid_sysid_translator_avalon_anti_slave_0_address;                                           // SysID_SysID_translator:av_address -> SysID:avs_SysID_address
	wire         sysid_sysid_translator_avalon_anti_slave_0_read;                                              // SysID_SysID_translator:av_read -> SysID:avs_SysID_read
	wire  [31:0] sysid_sysid_translator_avalon_anti_slave_0_readdata;                                          // SysID:avs_SysID_readdata -> SysID_SysID_translator:av_readdata
	wire         test_regwaitrw32_0_test_translator_avalon_anti_slave_0_waitrequest;                           // test_RegWaitRW32_0:avs_test_waitrequest -> test_RegWaitRW32_0_test_translator:av_waitrequest
	wire  [31:0] test_regwaitrw32_0_test_translator_avalon_anti_slave_0_writedata;                             // test_RegWaitRW32_0_test_translator:av_writedata -> test_RegWaitRW32_0:avs_test_writedata
	wire   [5:0] test_regwaitrw32_0_test_translator_avalon_anti_slave_0_address;                               // test_RegWaitRW32_0_test_translator:av_address -> test_RegWaitRW32_0:avs_test_address
	wire         test_regwaitrw32_0_test_translator_avalon_anti_slave_0_write;                                 // test_RegWaitRW32_0_test_translator:av_write -> test_RegWaitRW32_0:avs_test_write
	wire         test_regwaitrw32_0_test_translator_avalon_anti_slave_0_read;                                  // test_RegWaitRW32_0_test_translator:av_read -> test_RegWaitRW32_0:avs_test_read
	wire  [31:0] test_regwaitrw32_0_test_translator_avalon_anti_slave_0_readdata;                              // test_RegWaitRW32_0:avs_test_readdata -> test_RegWaitRW32_0_test_translator:av_readdata
	wire         test_regwaitrw32_0_test_translator_avalon_anti_slave_0_readdatavalid;                         // test_RegWaitRW32_0:avs_test_readdatavalid -> test_RegWaitRW32_0_test_translator:av_readdatavalid
	wire   [3:0] test_regwaitrw32_0_test_translator_avalon_anti_slave_0_byteenable;                            // test_RegWaitRW32_0_test_translator:av_byteenable -> test_RegWaitRW32_0:avs_test_byteenable
	wire         hps_tabby_m1_translator_avalon_universal_master_0_waitrequest;                                // HPS_Tabby_M1_translator_avalon_universal_master_0_agent:av_waitrequest -> HPS_Tabby_M1_translator:uav_waitrequest
	wire   [2:0] hps_tabby_m1_translator_avalon_universal_master_0_burstcount;                                 // HPS_Tabby_M1_translator:uav_burstcount -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] hps_tabby_m1_translator_avalon_universal_master_0_writedata;                                  // HPS_Tabby_M1_translator:uav_writedata -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] hps_tabby_m1_translator_avalon_universal_master_0_address;                                    // HPS_Tabby_M1_translator:uav_address -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:av_address
	wire         hps_tabby_m1_translator_avalon_universal_master_0_lock;                                       // HPS_Tabby_M1_translator:uav_lock -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:av_lock
	wire         hps_tabby_m1_translator_avalon_universal_master_0_write;                                      // HPS_Tabby_M1_translator:uav_write -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:av_write
	wire         hps_tabby_m1_translator_avalon_universal_master_0_read;                                       // HPS_Tabby_M1_translator:uav_read -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] hps_tabby_m1_translator_avalon_universal_master_0_readdata;                                   // HPS_Tabby_M1_translator_avalon_universal_master_0_agent:av_readdata -> HPS_Tabby_M1_translator:uav_readdata
	wire         hps_tabby_m1_translator_avalon_universal_master_0_debugaccess;                                // HPS_Tabby_M1_translator:uav_debugaccess -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] hps_tabby_m1_translator_avalon_universal_master_0_byteenable;                                 // HPS_Tabby_M1_translator:uav_byteenable -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:av_byteenable
	wire         hps_tabby_m1_translator_avalon_universal_master_0_readdatavalid;                              // HPS_Tabby_M1_translator_avalon_universal_master_0_agent:av_readdatavalid -> HPS_Tabby_M1_translator:uav_readdatavalid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // SysID_SysID_translator:uav_waitrequest -> SysID_SysID_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_burstcount -> SysID_SysID_translator:uav_burstcount
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_writedata;                           // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_writedata -> SysID_SysID_translator:uav_writedata
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_address;                             // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_address -> SysID_SysID_translator:uav_address
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_write;                               // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_write -> SysID_SysID_translator:uav_write
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_lock;                                // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_lock -> SysID_SysID_translator:uav_lock
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_read;                                // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_read -> SysID_SysID_translator:uav_read
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdata;                            // SysID_SysID_translator:uav_readdata -> SysID_SysID_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // SysID_SysID_translator:uav_readdatavalid -> SysID_SysID_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SysID_SysID_translator:uav_debugaccess
	wire   [3:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_byteenable -> SysID_SysID_translator:uav_byteenable
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [83:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_data;                         // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_data -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [83:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // test_RegWaitRW32_0_test_translator:uav_waitrequest -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_burstcount;              // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:m0_burstcount -> test_RegWaitRW32_0_test_translator:uav_burstcount
	wire  [31:0] test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_writedata;               // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:m0_writedata -> test_RegWaitRW32_0_test_translator:uav_writedata
	wire  [31:0] test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_address;                 // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:m0_address -> test_RegWaitRW32_0_test_translator:uav_address
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_write;                   // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:m0_write -> test_RegWaitRW32_0_test_translator:uav_write
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_lock;                    // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:m0_lock -> test_RegWaitRW32_0_test_translator:uav_lock
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_read;                    // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:m0_read -> test_RegWaitRW32_0_test_translator:uav_read
	wire  [31:0] test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdata;                // test_RegWaitRW32_0_test_translator:uav_readdata -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // test_RegWaitRW32_0_test_translator:uav_readdatavalid -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:m0_debugaccess -> test_RegWaitRW32_0_test_translator:uav_debugaccess
	wire   [3:0] test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_byteenable;              // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:m0_byteenable -> test_RegWaitRW32_0_test_translator:uav_byteenable
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_valid;            // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rf_source_valid -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [83:0] test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_data;             // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rf_source_data -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_ready;            // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [83:0] test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rf_sink_ready -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // HPS_Tabby_M1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_valid;                             // HPS_Tabby_M1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // HPS_Tabby_M1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [82:0] hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_data;                              // HPS_Tabby_M1_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router:sink_ready -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:cp_ready
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_valid;                               // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [82:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rp_data;                                // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router:sink_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent:rp_ready
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_valid;                   // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [82:0] test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_data;                    // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_001:sink_ready -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                  // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                        // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [82:0] addr_router_src_data;                                                                         // addr_router:src_data -> limiter:cmd_sink_data
	wire   [1:0] addr_router_src_channel;                                                                      // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                        // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                  // limiter:rsp_src_endofpacket -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                        // limiter:rsp_src_valid -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                // limiter:rsp_src_startofpacket -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [82:0] limiter_rsp_src_data;                                                                         // limiter:rsp_src_data -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] limiter_rsp_src_channel;                                                                      // limiter:rsp_src_channel -> HPS_Tabby_M1_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                        // HPS_Tabby_M1_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         cmd_xbar_demux_src0_endofpacket;                                                              // cmd_xbar_demux:src0_endofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                    // cmd_xbar_demux:src0_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                            // cmd_xbar_demux:src0_startofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [82:0] cmd_xbar_demux_src0_data;                                                                     // cmd_xbar_demux:src0_data -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_demux_src0_channel;                                                                  // cmd_xbar_demux:src0_channel -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src1_endofpacket;                                                              // cmd_xbar_demux:src1_endofpacket -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                    // cmd_xbar_demux:src1_valid -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                            // cmd_xbar_demux:src1_startofpacket -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [82:0] cmd_xbar_demux_src1_data;                                                                     // cmd_xbar_demux:src1_data -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_demux_src1_channel;                                                                  // cmd_xbar_demux:src1_channel -> test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                              // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                    // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                            // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [82:0] rsp_xbar_demux_src0_data;                                                                     // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [1:0] rsp_xbar_demux_src0_channel;                                                                  // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                    // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                          // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                        // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [82:0] rsp_xbar_demux_001_src0_data;                                                                 // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [1:0] rsp_xbar_demux_001_src0_channel;                                                              // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                  // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [82:0] limiter_cmd_src_data;                                                                         // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [1:0] limiter_cmd_src_channel;                                                                      // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                        // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                 // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                       // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                               // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [82:0] rsp_xbar_mux_src_data;                                                                        // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [1:0] rsp_xbar_mux_src_channel;                                                                     // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                       // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         cmd_xbar_demux_src0_ready;                                                                    // SysID_SysID_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire         id_router_src_endofpacket;                                                                    // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                          // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                  // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [82:0] id_router_src_data;                                                                           // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [1:0] id_router_src_channel;                                                                        // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                          // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_demux_src1_ready;                                                                    // test_RegWaitRW32_0_test_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire         id_router_001_src_endofpacket;                                                                // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                      // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                              // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [82:0] id_router_001_src_data;                                                                       // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [1:0] id_router_001_src_channel;                                                                    // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                      // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire   [1:0] limiter_cmd_valid_data;                                                                       // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [9:0] hps_tabby_events_irq;                                                                         // irq_synchronizer:sender_irq -> HPS_Tabby:inr_EVENTS_irq
	wire   [9:0] irq_synchronizer_receiver_irq;                                                                // irq_mapper:sender_irq -> irq_synchronizer:receiver_irq

	hps_tabby hps_tabby (
		.rso_MRST_reset       (hps_tabby_mrst_reset),       //   MRST.reset
		.cso_MCLK_clk         (hps_tabby_mclk_clk),         //   MCLK.clk
		.cso_H1CLK_clk        (),                           //  H1CLK.clk
		.cso_H2CLK_clk        (),                           //  H2CLK.clk
		.avm_M1_writedata     (hps_tabby_m1_writedata),     //     M1.writedata
		.avm_M1_readdata      (hps_tabby_m1_readdata),      //       .readdata
		.avm_M1_address       (hps_tabby_m1_address),       //       .address
		.avm_M1_byteenable    (hps_tabby_m1_byteenable),    //       .byteenable
		.avm_M1_write         (hps_tabby_m1_write),         //       .write
		.avm_M1_read          (hps_tabby_m1_read),          //       .read
		.avm_M1_begintransfer (hps_tabby_m1_begintransfer), //       .begintransfer
		.avm_M1_readdatavalid (hps_tabby_m1_readdatavalid), //       .readdatavalid
		.avm_M1_waitrequest   (hps_tabby_m1_waitrequest),   //       .waitrequest
		.inr_EVENTS_irq       (hps_tabby_events_irq),       // EVENTS.irq
		.coe_M1_RSTN          (m1_RSTN),                    // EXPORT.export
		.coe_M1_CLK           (m1_CLK),                     //       .export
		.coe_M1_ADDR          (m1_ADDR),                    //       .export
		.coe_M1_DATA          (m1_DATA),                    //       .export
		.coe_M1_CSN           (m1_CSN),                     //       .export
		.coe_M1_BEN           (m1_BEN),                     //       .export
		.coe_M1_RDN           (m1_RDN),                     //       .export
		.coe_M1_WRN           (m1_WRN),                     //       .export
		.coe_M1_WAITN         (m1_WAITN),                   //       .export
		.coe_M1_EINT          (m1_EINT)                     //       .export
	);

	basic_SysID sysid (
		.rsi_MRST_reset        (hps_tabby_mrst_reset),                                   //  MRST.reset
		.csi_MCLK_clk          (hps_tabby_mclk_clk),                                     //  MCLK.clk
		.avs_SysID_readdata    (sysid_sysid_translator_avalon_anti_slave_0_readdata),    // SysID.readdata
		.avs_SysID_address     (sysid_sysid_translator_avalon_anti_slave_0_address),     //      .address
		.avs_SysID_read        (sysid_sysid_translator_avalon_anti_slave_0_read),        //      .read
		.avs_SysID_waitrequest (sysid_sysid_translator_avalon_anti_slave_0_waitrequest)  //      .waitrequest
	);

	test_RegWaitRW32 test_regwaitrw32_0 (
		.rsi_MRST_reset         (hps_tabby_mrst_reset),                                                 // MRST.reset
		.csi_MCLK_clk           (hps_tabby_mclk_clk),                                                   // MCLK.clk
		.avs_test_writedata     (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_writedata),     // test.writedata
		.avs_test_readdata      (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_readdata),      //     .readdata
		.avs_test_address       (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_address),       //     .address
		.avs_test_byteenable    (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_byteenable),    //     .byteenable
		.avs_test_write         (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_write),         //     .write
		.avs_test_read          (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_read),          //     .read
		.avs_test_waitrequest   (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_waitrequest),   //     .waitrequest
		.avs_test_readdatavalid (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_readdatavalid)  //     .readdatavalid
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (30),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (1),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (0),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) hps_tabby_m1_translator (
		.clk                   (hps_tabby_mclk_clk),                                              //                       clk.clk
		.reset                 (hps_tabby_mrst_reset),                                            //                     reset.reset
		.uav_address           (hps_tabby_m1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (hps_tabby_m1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (hps_tabby_m1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (hps_tabby_m1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (hps_tabby_m1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (hps_tabby_m1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (hps_tabby_m1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (hps_tabby_m1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (hps_tabby_m1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (hps_tabby_m1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (hps_tabby_m1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (hps_tabby_m1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (hps_tabby_m1_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (hps_tabby_m1_byteenable),                                         //                          .byteenable
		.av_begintransfer      (hps_tabby_m1_begintransfer),                                      //                          .begintransfer
		.av_read               (hps_tabby_m1_read),                                               //                          .read
		.av_readdata           (hps_tabby_m1_readdata),                                           //                          .readdata
		.av_readdatavalid      (hps_tabby_m1_readdatavalid),                                      //                          .readdatavalid
		.av_write              (hps_tabby_m1_write),                                              //                          .write
		.av_writedata          (hps_tabby_m1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                            //               (terminated)
		.av_chipselect         (1'b0),                                                            //               (terminated)
		.av_lock               (1'b0),                                                            //               (terminated)
		.av_debugaccess        (1'b0),                                                            //               (terminated)
		.uav_clken             (),                                                                //               (terminated)
		.av_clken              (1'b1)                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_sysid_translator (
		.clk                   (hps_tabby_mclk_clk),                                                     //                      clk.clk
		.reset                 (hps_tabby_mrst_reset),                                                   //                    reset.reset
		.uav_address           (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_sysid_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_read               (sysid_sysid_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sysid_sysid_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (sysid_sysid_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_write              (),                                                                       //              (terminated)
		.av_writedata          (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_chipselect         (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (6),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) test_regwaitrw32_0_test_translator (
		.clk                   (hps_tabby_mclk_clk),                                                                 //                      clk.clk
		.reset                 (hps_tabby_mrst_reset),                                                               //                    reset.reset
		.uav_address           (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (test_regwaitrw32_0_test_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_chipselect         (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (82),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (81),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7)
	) hps_tabby_m1_translator_avalon_universal_master_0_agent (
		.clk              (hps_tabby_mclk_clk),                                                       //       clk.clk
		.reset            (hps_tabby_mrst_reset),                                                     // clk_reset.reset
		.av_address       (hps_tabby_m1_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (hps_tabby_m1_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (hps_tabby_m1_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (hps_tabby_m1_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (hps_tabby_m1_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (hps_tabby_m1_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (hps_tabby_m1_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (hps_tabby_m1_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (hps_tabby_m1_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (hps_tabby_m1_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (hps_tabby_m1_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                    //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                     //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                  //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                     //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (82),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_sysid_translator_avalon_universal_slave_0_agent (
		.clk                     (hps_tabby_mclk_clk),                                                               //             clk.clk
		.reset                   (hps_tabby_mrst_reset),                                                             //       clk_reset.reset
		.m0_address              (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                      //                .channel
		.rf_sink_ready           (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (hps_tabby_mclk_clk),                                                               //       clk.clk
		.reset             (hps_tabby_mrst_reset),                                                             // clk_reset.reset
		.in_data           (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (82),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent (
		.clk                     (hps_tabby_mclk_clk),                                                                           //             clk.clk
		.reset                   (hps_tabby_mrst_reset),                                                                         //       clk_reset.reset
		.m0_address              (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                                  //                .channel
		.rf_sink_ready           (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (hps_tabby_mclk_clk),                                                                           //       clk.clk
		.reset             (hps_tabby_mrst_reset),                                                                         // clk_reset.reset
		.in_data           (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	frontier_addr_router addr_router (
		.sink_ready         (hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hps_tabby_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (hps_tabby_mclk_clk),                                                       //       clk.clk
		.reset              (hps_tabby_mrst_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_src_valid),                                                    //          .valid
		.src_data           (addr_router_src_data),                                                     //          .data
		.src_channel        (addr_router_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                               //          .endofpacket
	);

	frontier_id_router id_router (
		.sink_ready         (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (hps_tabby_mclk_clk),                                                     //       clk.clk
		.reset              (hps_tabby_mrst_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                    //       src.ready
		.src_valid          (id_router_src_valid),                                                    //          .valid
		.src_data           (id_router_src_data),                                                     //          .data
		.src_channel        (id_router_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                               //          .endofpacket
	);

	frontier_id_router id_router_001 (
		.sink_ready         (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (test_regwaitrw32_0_test_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (hps_tabby_mclk_clk),                                                                 //       clk.clk
		.reset              (hps_tabby_mrst_reset),                                                               // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                            //       src.ready
		.src_valid          (id_router_001_src_valid),                                                            //          .valid
		.src_data           (id_router_001_src_data),                                                             //          .data
		.src_channel        (id_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (81),
		.PKT_DEST_ID_L             (81),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (2),
		.VALID_WIDTH               (2),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (hps_tabby_mclk_clk),             //       clk.clk
		.reset                  (hps_tabby_mrst_reset),           // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	frontier_cmd_xbar_demux cmd_xbar_demux (
		.clk                (hps_tabby_mclk_clk),                //        clk.clk
		.reset              (hps_tabby_mrst_reset),              //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //           .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux (
		.clk                (hps_tabby_mclk_clk),                //       clk.clk
		.reset              (hps_tabby_mrst_reset),              // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (hps_tabby_mclk_clk),                    //       clk.clk
		.reset              (hps_tabby_mrst_reset),                  // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (hps_tabby_mclk_clk),                    //       clk.clk
		.reset               (hps_tabby_mrst_reset),                  // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	frontier_irq_mapper irq_mapper (
		.clk        (hps_tabby_mclk_clk),            //       clk.clk
		.reset      (hps_tabby_mrst_reset),          // clk_reset.reset
		.sender_irq (irq_synchronizer_receiver_irq)  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (10)
	) irq_synchronizer (
		.receiver_clk   (hps_tabby_mclk_clk),            //       receiver_clk.clk
		.sender_clk     (hps_tabby_mclk_clk),            //         sender_clk.clk
		.receiver_reset (hps_tabby_mrst_reset),          // receiver_clk_reset.reset
		.sender_reset   (hps_tabby_mrst_reset),          //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq), //           receiver.irq
		.sender_irq     (hps_tabby_events_irq)           //             sender.irq
	);

endmodule
