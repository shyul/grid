// frontier.v

// Generated using ACDS version 11.1sp2 259 at 2012.07.20.17:04:57

`timescale 1 ps / 1 ps
module frontier (
		output wire        led_f3_R,       // led_f3.R
		output wire        led_f3_G,       //       .G
		output wire        led_f3_B,       //       .B
		output wire        led_f2_R,       // led_f2.R
		output wire        led_f2_G,       //       .G
		output wire        led_f2_B,       //       .B
		inout  wire        slot_a_P0,      // slot_a.P0
		inout  wire        slot_a_P1,      //       .P1
		inout  wire        slot_a_P2,      //       .P2
		inout  wire        slot_a_P3,      //       .P3
		inout  wire        slot_a_P4,      //       .P4
		inout  wire        slot_a_P5,      //       .P5
		inout  wire        slot_a_P6,      //       .P6
		inout  wire        slot_a_P7,      //       .P7
		inout  wire        slot_a_P8,      //       .P8
		inout  wire        slot_a_P9,      //       .P9
		inout  wire        slot_a_P10,     //       .P10
		inout  wire        slot_a_P11,     //       .P11
		inout  wire        slot_a_P12,     //       .P12
		inout  wire        slot_a_P13,     //       .P13
		inout  wire        slot_a_P14,     //       .P14
		inout  wire        slot_a_P15,     //       .P15
		inout  wire        slot_a_P16,     //       .P16
		inout  wire        slot_a_P17,     //       .P17
		inout  wire        slot_a_P18,     //       .P18
		inout  wire        slot_a_P19,     //       .P19
		inout  wire        slot_a_P20,     //       .P20
		inout  wire        slot_a_P21,     //       .P21
		inout  wire        slot_a_P22,     //       .P22
		inout  wire        slot_a_P23,     //       .P23
		inout  wire        slot_a_P24,     //       .P24
		inout  wire        slot_a_P25,     //       .P25
		inout  wire        slot_b_P0,      // slot_b.P0
		inout  wire        slot_b_P1,      //       .P1
		inout  wire        slot_b_P2,      //       .P2
		inout  wire        slot_b_P3,      //       .P3
		inout  wire        slot_b_P4,      //       .P4
		inout  wire        slot_b_P5,      //       .P5
		inout  wire        slot_b_P6,      //       .P6
		inout  wire        slot_b_P7,      //       .P7
		inout  wire        slot_b_P8,      //       .P8
		inout  wire        slot_b_P9,      //       .P9
		inout  wire        slot_b_P10,     //       .P10
		inout  wire        slot_b_P11,     //       .P11
		inout  wire        slot_b_P12,     //       .P12
		inout  wire        slot_b_P13,     //       .P13
		inout  wire        slot_b_P14,     //       .P14
		inout  wire        slot_b_P15,     //       .P15
		inout  wire        slot_b_P16,     //       .P16
		inout  wire        slot_b_P17,     //       .P17
		inout  wire        slot_b_P18,     //       .P18
		inout  wire        slot_b_P19,     //       .P19
		inout  wire        slot_b_P20,     //       .P20
		inout  wire        slot_b_P21,     //       .P21
		inout  wire        slot_b_P22,     //       .P22
		inout  wire        slot_b_P23,     //       .P23
		inout  wire        slot_b_P24,     //       .P24
		inout  wire        slot_b_P25,     //       .P25
		input  wire        m1_RSTN,        //     m1.RSTN
		input  wire        m1_CLK,         //       .CLK
		input  wire [21:0] m1_ADDR,        //       .ADDR
		inout  wire [31:0] m1_DATA,        //       .DATA
		input  wire [3:0]  m1_CSN,         //       .CSN
		input  wire [3:0]  m1_BEN,         //       .BEN
		input  wire        m1_RDN,         //       .RDN
		input  wire        m1_WRN,         //       .WRN
		output wire        m1_WAITN,       //       .WAITN
		output wire [9:0]  m1_EINT,        //       .EINT
		output wire        led_f0_R,       // led_f0.R
		output wire        led_f0_G,       //       .G
		output wire        led_f0_B,       //       .B
		output wire        led_f1_R,       // led_f1.R
		output wire        led_f1_G,       //       .G
		output wire        led_f1_B,       //       .B
		input  wire        shield_A_OCN,   // shield.A_OCN
		output wire        shield_A_PWREN, //       .A_PWREN
		output wire        shield_A_HOE,   //       .A_HOE
		output wire        shield_A_LOE,   //       .A_LOE
		input  wire        shield_B_OCN,   //       .B_OCN
		output wire        shield_B_PWREN, //       .B_PWREN
		output wire        shield_B_HOE,   //       .B_HOE
		output wire        shield_B_LOE    //       .B_LOE
	);

	wire         sam9_mrst_reset;                                                                        // SAM9:rso_MRST_reset -> [FuncLED_0:rsi_MRST_reset, FuncLED_0_LEDD_translator:reset, FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:reset, FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FuncLED_1:rsi_MRST_reset, FuncLED_1_LEDD_translator:reset, FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:reset, FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FuncLED_2:rsi_MRST_reset, FuncLED_2_LEDD_translator:reset, FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:reset, FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FuncLED_3:rsi_MRST_reset, FuncLED_3_LEDD_translator:reset, FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:reset, FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SAM9_M1_translator:reset, SAM9_M1_translator_avalon_universal_master_0_agent:reset, Shield_Admin:rsi_MRST_reset, Shield_Admin_Ctrl_translator:reset, Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:reset, Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shield_PIO_A:rsi_MRST_reset, Shield_PIO_A_gpio_translator:reset, Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:reset, Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Shield_PIO_B:rsi_MRST_reset, Shield_PIO_B_gpio_translator:reset, Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:reset, Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SysID:rsi_MRST_reset, SysID_SysID_translator:reset, SysID_SysID_translator_avalon_universal_slave_0_agent:reset, SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, cmd_xbar_demux:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, irq_mapper:reset, irq_synchronizer:receiver_reset, irq_synchronizer:sender_reset, limiter:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_mux:reset, test_LEDState_0:rsi_MRST_reset, test_LEDState_1:rsi_MRST_reset, test_LEDState_2:rsi_MRST_reset, test_LEDState_3:rsi_MRST_reset]
	wire         sam9_mclk_clk;                                                                          // SAM9:cso_MCLK_clk -> [FuncLED_0:csi_MCLK_clk, FuncLED_0_LEDD_translator:clk, FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:clk, FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, FuncLED_1:csi_MCLK_clk, FuncLED_1_LEDD_translator:clk, FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:clk, FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, FuncLED_2:csi_MCLK_clk, FuncLED_2_LEDD_translator:clk, FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:clk, FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, FuncLED_3:csi_MCLK_clk, FuncLED_3_LEDD_translator:clk, FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:clk, FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, SAM9_M1_translator:clk, SAM9_M1_translator_avalon_universal_master_0_agent:clk, Shield_Admin:csi_MCLK_clk, Shield_Admin_Ctrl_translator:clk, Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:clk, Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shield_PIO_A:csi_MCLK_clk, Shield_PIO_A_gpio_translator:clk, Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:clk, Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, Shield_PIO_B:csi_MCLK_clk, Shield_PIO_B_gpio_translator:clk, Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:clk, Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, SysID:csi_MCLK_clk, SysID_SysID_translator:clk, SysID_SysID_translator_avalon_universal_slave_0_agent:clk, SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, cmd_xbar_demux:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, irq_mapper:clk, irq_synchronizer:receiver_clk, irq_synchronizer:sender_clk, limiter:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_mux:clk, test_LEDState_0:csi_MCLK_clk, test_LEDState_1:csi_MCLK_clk, test_LEDState_2:csi_MCLK_clk, test_LEDState_3:csi_MCLK_clk]
	wire         test_ledstate_1_leds_valid;                                                             // test_LEDState_1:aso_LEDS_valid -> FuncLED_1:asi_LEDS_valid
	wire  [23:0] test_ledstate_1_leds_data;                                                              // test_LEDState_1:aso_LEDS_data -> FuncLED_1:asi_LEDS_data
	wire         test_ledstate_1_leds_ready;                                                             // FuncLED_1:asi_LEDS_ready -> test_LEDState_1:aso_LEDS_ready
	wire         test_ledstate_2_leds_valid;                                                             // test_LEDState_2:aso_LEDS_valid -> FuncLED_2:asi_LEDS_valid
	wire  [23:0] test_ledstate_2_leds_data;                                                              // test_LEDState_2:aso_LEDS_data -> FuncLED_2:asi_LEDS_data
	wire         test_ledstate_2_leds_ready;                                                             // FuncLED_2:asi_LEDS_ready -> test_LEDState_2:aso_LEDS_ready
	wire         test_ledstate_3_leds_valid;                                                             // test_LEDState_3:aso_LEDS_valid -> FuncLED_3:asi_LEDS_valid
	wire  [23:0] test_ledstate_3_leds_data;                                                              // test_LEDState_3:aso_LEDS_data -> FuncLED_3:asi_LEDS_data
	wire         test_ledstate_3_leds_ready;                                                             // FuncLED_3:asi_LEDS_ready -> test_LEDState_3:aso_LEDS_ready
	wire         test_ledstate_0_leds_valid;                                                             // test_LEDState_0:aso_LEDS_valid -> FuncLED_0:asi_LEDS_valid
	wire  [23:0] test_ledstate_0_leds_data;                                                              // test_LEDState_0:aso_LEDS_data -> FuncLED_0:asi_LEDS_data
	wire         test_ledstate_0_leds_ready;                                                             // FuncLED_0:asi_LEDS_ready -> test_LEDState_0:aso_LEDS_ready
	wire         sam9_m1_waitrequest;                                                                    // SAM9_M1_translator:av_waitrequest -> SAM9:avm_M1_waitrequest
	wire  [31:0] sam9_m1_address;                                                                        // SAM9:avm_M1_address -> SAM9_M1_translator:av_address
	wire  [31:0] sam9_m1_writedata;                                                                      // SAM9:avm_M1_writedata -> SAM9_M1_translator:av_writedata
	wire         sam9_m1_write;                                                                          // SAM9:avm_M1_write -> SAM9_M1_translator:av_write
	wire         sam9_m1_read;                                                                           // SAM9:avm_M1_read -> SAM9_M1_translator:av_read
	wire  [31:0] sam9_m1_readdata;                                                                       // SAM9_M1_translator:av_readdata -> SAM9:avm_M1_readdata
	wire         sam9_m1_begintransfer;                                                                  // SAM9:avm_M1_begintransfer -> SAM9_M1_translator:av_begintransfer
	wire         sam9_m1_readdatavalid;                                                                  // SAM9_M1_translator:av_readdatavalid -> SAM9:avm_M1_readdatavalid
	wire   [3:0] sam9_m1_byteenable;                                                                     // SAM9:avm_M1_byteenable -> SAM9_M1_translator:av_byteenable
	wire         sysid_sysid_translator_avalon_anti_slave_0_waitrequest;                                 // SysID:avs_SysID_waitrequest -> SysID_SysID_translator:av_waitrequest
	wire         sysid_sysid_translator_avalon_anti_slave_0_read;                                        // SysID_SysID_translator:av_read -> SysID:avs_SysID_read
	wire  [31:0] sysid_sysid_translator_avalon_anti_slave_0_readdata;                                    // SysID:avs_SysID_readdata -> SysID_SysID_translator:av_readdata
	wire         funcled_0_ledd_translator_avalon_anti_slave_0_waitrequest;                              // FuncLED_0:avs_LEDD_waitrequest -> FuncLED_0_LEDD_translator:av_waitrequest
	wire  [31:0] funcled_0_ledd_translator_avalon_anti_slave_0_writedata;                                // FuncLED_0_LEDD_translator:av_writedata -> FuncLED_0:avs_LEDD_writedata
	wire         funcled_0_ledd_translator_avalon_anti_slave_0_write;                                    // FuncLED_0_LEDD_translator:av_write -> FuncLED_0:avs_LEDD_write
	wire         funcled_0_ledd_translator_avalon_anti_slave_0_read;                                     // FuncLED_0_LEDD_translator:av_read -> FuncLED_0:avs_LEDD_read
	wire  [31:0] funcled_0_ledd_translator_avalon_anti_slave_0_readdata;                                 // FuncLED_0:avs_LEDD_readdata -> FuncLED_0_LEDD_translator:av_readdata
	wire   [3:0] funcled_0_ledd_translator_avalon_anti_slave_0_byteenable;                               // FuncLED_0_LEDD_translator:av_byteenable -> FuncLED_0:avs_LEDD_byteenable
	wire         funcled_1_ledd_translator_avalon_anti_slave_0_waitrequest;                              // FuncLED_1:avs_LEDD_waitrequest -> FuncLED_1_LEDD_translator:av_waitrequest
	wire  [31:0] funcled_1_ledd_translator_avalon_anti_slave_0_writedata;                                // FuncLED_1_LEDD_translator:av_writedata -> FuncLED_1:avs_LEDD_writedata
	wire         funcled_1_ledd_translator_avalon_anti_slave_0_write;                                    // FuncLED_1_LEDD_translator:av_write -> FuncLED_1:avs_LEDD_write
	wire         funcled_1_ledd_translator_avalon_anti_slave_0_read;                                     // FuncLED_1_LEDD_translator:av_read -> FuncLED_1:avs_LEDD_read
	wire  [31:0] funcled_1_ledd_translator_avalon_anti_slave_0_readdata;                                 // FuncLED_1:avs_LEDD_readdata -> FuncLED_1_LEDD_translator:av_readdata
	wire   [3:0] funcled_1_ledd_translator_avalon_anti_slave_0_byteenable;                               // FuncLED_1_LEDD_translator:av_byteenable -> FuncLED_1:avs_LEDD_byteenable
	wire         funcled_2_ledd_translator_avalon_anti_slave_0_waitrequest;                              // FuncLED_2:avs_LEDD_waitrequest -> FuncLED_2_LEDD_translator:av_waitrequest
	wire  [31:0] funcled_2_ledd_translator_avalon_anti_slave_0_writedata;                                // FuncLED_2_LEDD_translator:av_writedata -> FuncLED_2:avs_LEDD_writedata
	wire         funcled_2_ledd_translator_avalon_anti_slave_0_write;                                    // FuncLED_2_LEDD_translator:av_write -> FuncLED_2:avs_LEDD_write
	wire         funcled_2_ledd_translator_avalon_anti_slave_0_read;                                     // FuncLED_2_LEDD_translator:av_read -> FuncLED_2:avs_LEDD_read
	wire  [31:0] funcled_2_ledd_translator_avalon_anti_slave_0_readdata;                                 // FuncLED_2:avs_LEDD_readdata -> FuncLED_2_LEDD_translator:av_readdata
	wire   [3:0] funcled_2_ledd_translator_avalon_anti_slave_0_byteenable;                               // FuncLED_2_LEDD_translator:av_byteenable -> FuncLED_2:avs_LEDD_byteenable
	wire         funcled_3_ledd_translator_avalon_anti_slave_0_waitrequest;                              // FuncLED_3:avs_LEDD_waitrequest -> FuncLED_3_LEDD_translator:av_waitrequest
	wire  [31:0] funcled_3_ledd_translator_avalon_anti_slave_0_writedata;                                // FuncLED_3_LEDD_translator:av_writedata -> FuncLED_3:avs_LEDD_writedata
	wire         funcled_3_ledd_translator_avalon_anti_slave_0_write;                                    // FuncLED_3_LEDD_translator:av_write -> FuncLED_3:avs_LEDD_write
	wire         funcled_3_ledd_translator_avalon_anti_slave_0_read;                                     // FuncLED_3_LEDD_translator:av_read -> FuncLED_3:avs_LEDD_read
	wire  [31:0] funcled_3_ledd_translator_avalon_anti_slave_0_readdata;                                 // FuncLED_3:avs_LEDD_readdata -> FuncLED_3_LEDD_translator:av_readdata
	wire   [3:0] funcled_3_ledd_translator_avalon_anti_slave_0_byteenable;                               // FuncLED_3_LEDD_translator:av_byteenable -> FuncLED_3:avs_LEDD_byteenable
	wire         shield_admin_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // Shield_Admin:avs_Ctrl_waitrequest -> Shield_Admin_Ctrl_translator:av_waitrequest
	wire  [31:0] shield_admin_ctrl_translator_avalon_anti_slave_0_writedata;                             // Shield_Admin_Ctrl_translator:av_writedata -> Shield_Admin:avs_Ctrl_writedata
	wire         shield_admin_ctrl_translator_avalon_anti_slave_0_write;                                 // Shield_Admin_Ctrl_translator:av_write -> Shield_Admin:avs_Ctrl_write
	wire         shield_admin_ctrl_translator_avalon_anti_slave_0_read;                                  // Shield_Admin_Ctrl_translator:av_read -> Shield_Admin:avs_Ctrl_read
	wire  [31:0] shield_admin_ctrl_translator_avalon_anti_slave_0_readdata;                              // Shield_Admin:avs_Ctrl_readdata -> Shield_Admin_Ctrl_translator:av_readdata
	wire   [3:0] shield_admin_ctrl_translator_avalon_anti_slave_0_byteenable;                            // Shield_Admin_Ctrl_translator:av_byteenable -> Shield_Admin:avs_Ctrl_byteenable
	wire         shield_pio_a_gpio_translator_avalon_anti_slave_0_waitrequest;                           // Shield_PIO_A:avs_gpio_waitrequest -> Shield_PIO_A_gpio_translator:av_waitrequest
	wire  [31:0] shield_pio_a_gpio_translator_avalon_anti_slave_0_writedata;                             // Shield_PIO_A_gpio_translator:av_writedata -> Shield_PIO_A:avs_gpio_writedata
	wire   [4:0] shield_pio_a_gpio_translator_avalon_anti_slave_0_address;                               // Shield_PIO_A_gpio_translator:av_address -> Shield_PIO_A:avs_gpio_address
	wire         shield_pio_a_gpio_translator_avalon_anti_slave_0_write;                                 // Shield_PIO_A_gpio_translator:av_write -> Shield_PIO_A:avs_gpio_write
	wire         shield_pio_a_gpio_translator_avalon_anti_slave_0_read;                                  // Shield_PIO_A_gpio_translator:av_read -> Shield_PIO_A:avs_gpio_read
	wire  [31:0] shield_pio_a_gpio_translator_avalon_anti_slave_0_readdata;                              // Shield_PIO_A:avs_gpio_readdata -> Shield_PIO_A_gpio_translator:av_readdata
	wire   [3:0] shield_pio_a_gpio_translator_avalon_anti_slave_0_byteenable;                            // Shield_PIO_A_gpio_translator:av_byteenable -> Shield_PIO_A:avs_gpio_byteenable
	wire         shield_pio_b_gpio_translator_avalon_anti_slave_0_waitrequest;                           // Shield_PIO_B:avs_gpio_waitrequest -> Shield_PIO_B_gpio_translator:av_waitrequest
	wire  [31:0] shield_pio_b_gpio_translator_avalon_anti_slave_0_writedata;                             // Shield_PIO_B_gpio_translator:av_writedata -> Shield_PIO_B:avs_gpio_writedata
	wire   [4:0] shield_pio_b_gpio_translator_avalon_anti_slave_0_address;                               // Shield_PIO_B_gpio_translator:av_address -> Shield_PIO_B:avs_gpio_address
	wire         shield_pio_b_gpio_translator_avalon_anti_slave_0_write;                                 // Shield_PIO_B_gpio_translator:av_write -> Shield_PIO_B:avs_gpio_write
	wire         shield_pio_b_gpio_translator_avalon_anti_slave_0_read;                                  // Shield_PIO_B_gpio_translator:av_read -> Shield_PIO_B:avs_gpio_read
	wire  [31:0] shield_pio_b_gpio_translator_avalon_anti_slave_0_readdata;                              // Shield_PIO_B:avs_gpio_readdata -> Shield_PIO_B_gpio_translator:av_readdata
	wire   [3:0] shield_pio_b_gpio_translator_avalon_anti_slave_0_byteenable;                            // Shield_PIO_B_gpio_translator:av_byteenable -> Shield_PIO_B:avs_gpio_byteenable
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // FuncLED_0_LEDD_translator:uav_waitrequest -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> FuncLED_0_LEDD_translator:uav_burstcount
	wire  [31:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                  // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> FuncLED_0_LEDD_translator:uav_writedata
	wire  [31:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_address;                    // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> FuncLED_0_LEDD_translator:uav_address
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_write;                      // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> FuncLED_0_LEDD_translator:uav_write
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                       // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> FuncLED_0_LEDD_translator:uav_lock
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_read;                       // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> FuncLED_0_LEDD_translator:uav_read
	wire  [31:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                   // FuncLED_0_LEDD_translator:uav_readdata -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // FuncLED_0_LEDD_translator:uav_readdatavalid -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FuncLED_0_LEDD_translator:uav_debugaccess
	wire   [3:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> FuncLED_0_LEDD_translator:uav_byteenable
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;               // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;               // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // SysID_SysID_translator:uav_waitrequest -> SysID_SysID_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_burstcount -> SysID_SysID_translator:uav_burstcount
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_writedata;                     // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_writedata -> SysID_SysID_translator:uav_writedata
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_address;                       // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_address -> SysID_SysID_translator:uav_address
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_write;                         // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_write -> SysID_SysID_translator:uav_write
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_lock;                          // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_lock -> SysID_SysID_translator:uav_lock
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_read;                          // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_read -> SysID_SysID_translator:uav_read
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdata;                      // SysID_SysID_translator:uav_readdata -> SysID_SysID_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // SysID_SysID_translator:uav_readdatavalid -> SysID_SysID_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SysID_SysID_translator:uav_debugaccess
	wire   [3:0] sysid_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // SysID_SysID_translator_avalon_universal_slave_0_agent:m0_byteenable -> SysID_SysID_translator:uav_byteenable
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_data;                   // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_data -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // SysID_SysID_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sam9_m1_translator_avalon_universal_master_0_waitrequest;                               // SAM9_M1_translator_avalon_universal_master_0_agent:av_waitrequest -> SAM9_M1_translator:uav_waitrequest
	wire   [2:0] sam9_m1_translator_avalon_universal_master_0_burstcount;                                // SAM9_M1_translator:uav_burstcount -> SAM9_M1_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] sam9_m1_translator_avalon_universal_master_0_writedata;                                 // SAM9_M1_translator:uav_writedata -> SAM9_M1_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] sam9_m1_translator_avalon_universal_master_0_address;                                   // SAM9_M1_translator:uav_address -> SAM9_M1_translator_avalon_universal_master_0_agent:av_address
	wire         sam9_m1_translator_avalon_universal_master_0_lock;                                      // SAM9_M1_translator:uav_lock -> SAM9_M1_translator_avalon_universal_master_0_agent:av_lock
	wire         sam9_m1_translator_avalon_universal_master_0_write;                                     // SAM9_M1_translator:uav_write -> SAM9_M1_translator_avalon_universal_master_0_agent:av_write
	wire         sam9_m1_translator_avalon_universal_master_0_read;                                      // SAM9_M1_translator:uav_read -> SAM9_M1_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] sam9_m1_translator_avalon_universal_master_0_readdata;                                  // SAM9_M1_translator_avalon_universal_master_0_agent:av_readdata -> SAM9_M1_translator:uav_readdata
	wire         sam9_m1_translator_avalon_universal_master_0_debugaccess;                               // SAM9_M1_translator:uav_debugaccess -> SAM9_M1_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] sam9_m1_translator_avalon_universal_master_0_byteenable;                                // SAM9_M1_translator:uav_byteenable -> SAM9_M1_translator_avalon_universal_master_0_agent:av_byteenable
	wire         sam9_m1_translator_avalon_universal_master_0_readdatavalid;                             // SAM9_M1_translator_avalon_universal_master_0_agent:av_readdatavalid -> SAM9_M1_translator:uav_readdatavalid
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shield_PIO_A_gpio_translator:uav_waitrequest -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shield_PIO_A_gpio_translator:uav_burstcount
	wire  [31:0] shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:m0_writedata -> Shield_PIO_A_gpio_translator:uav_writedata
	wire  [31:0] shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_address;                 // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:m0_address -> Shield_PIO_A_gpio_translator:uav_address
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_write;                   // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:m0_write -> Shield_PIO_A_gpio_translator:uav_write
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:m0_lock -> Shield_PIO_A_gpio_translator:uav_lock
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_read;                    // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:m0_read -> Shield_PIO_A_gpio_translator:uav_read
	wire  [31:0] shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shield_PIO_A_gpio_translator:uav_readdata -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shield_PIO_A_gpio_translator:uav_readdatavalid -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shield_PIO_A_gpio_translator:uav_debugaccess
	wire   [3:0] shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shield_PIO_A_gpio_translator:uav_byteenable
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rf_source_data -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // FuncLED_3_LEDD_translator:uav_waitrequest -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> FuncLED_3_LEDD_translator:uav_burstcount
	wire  [31:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                  // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> FuncLED_3_LEDD_translator:uav_writedata
	wire  [31:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_address;                    // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> FuncLED_3_LEDD_translator:uav_address
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_write;                      // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> FuncLED_3_LEDD_translator:uav_write
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                       // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> FuncLED_3_LEDD_translator:uav_lock
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_read;                       // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> FuncLED_3_LEDD_translator:uav_read
	wire  [31:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                   // FuncLED_3_LEDD_translator:uav_readdata -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // FuncLED_3_LEDD_translator:uav_readdatavalid -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FuncLED_3_LEDD_translator:uav_debugaccess
	wire   [3:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> FuncLED_3_LEDD_translator:uav_byteenable
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;               // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;               // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shield_Admin_Ctrl_translator:uav_waitrequest -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shield_Admin_Ctrl_translator:uav_burstcount
	wire  [31:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> Shield_Admin_Ctrl_translator:uav_writedata
	wire  [31:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_address -> Shield_Admin_Ctrl_translator:uav_address
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_write -> Shield_Admin_Ctrl_translator:uav_write
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> Shield_Admin_Ctrl_translator:uav_lock
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_read -> Shield_Admin_Ctrl_translator:uav_read
	wire  [31:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shield_Admin_Ctrl_translator:uav_readdata -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shield_Admin_Ctrl_translator:uav_readdatavalid -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shield_Admin_Ctrl_translator:uav_debugaccess
	wire   [3:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shield_Admin_Ctrl_translator:uav_byteenable
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // FuncLED_2_LEDD_translator:uav_waitrequest -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> FuncLED_2_LEDD_translator:uav_burstcount
	wire  [31:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                  // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> FuncLED_2_LEDD_translator:uav_writedata
	wire  [31:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_address;                    // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> FuncLED_2_LEDD_translator:uav_address
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_write;                      // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> FuncLED_2_LEDD_translator:uav_write
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                       // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> FuncLED_2_LEDD_translator:uav_lock
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_read;                       // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> FuncLED_2_LEDD_translator:uav_read
	wire  [31:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                   // FuncLED_2_LEDD_translator:uav_readdata -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // FuncLED_2_LEDD_translator:uav_readdatavalid -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FuncLED_2_LEDD_translator:uav_debugaccess
	wire   [3:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> FuncLED_2_LEDD_translator:uav_byteenable
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;               // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;               // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // FuncLED_1_LEDD_translator:uav_waitrequest -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> FuncLED_1_LEDD_translator:uav_burstcount
	wire  [31:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                  // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> FuncLED_1_LEDD_translator:uav_writedata
	wire  [31:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_address;                    // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> FuncLED_1_LEDD_translator:uav_address
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_write;                      // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> FuncLED_1_LEDD_translator:uav_write
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                       // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> FuncLED_1_LEDD_translator:uav_lock
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_read;                       // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> FuncLED_1_LEDD_translator:uav_read
	wire  [31:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                   // FuncLED_1_LEDD_translator:uav_readdata -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // FuncLED_1_LEDD_translator:uav_readdatavalid -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FuncLED_1_LEDD_translator:uav_debugaccess
	wire   [3:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> FuncLED_1_LEDD_translator:uav_byteenable
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;               // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;               // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Shield_PIO_B_gpio_translator:uav_waitrequest -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:m0_burstcount -> Shield_PIO_B_gpio_translator:uav_burstcount
	wire  [31:0] shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_writedata;               // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:m0_writedata -> Shield_PIO_B_gpio_translator:uav_writedata
	wire  [31:0] shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_address;                 // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:m0_address -> Shield_PIO_B_gpio_translator:uav_address
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_write;                   // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:m0_write -> Shield_PIO_B_gpio_translator:uav_write
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_lock;                    // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:m0_lock -> Shield_PIO_B_gpio_translator:uav_lock
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_read;                    // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:m0_read -> Shield_PIO_B_gpio_translator:uav_read
	wire  [31:0] shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_readdata;                // Shield_PIO_B_gpio_translator:uav_readdata -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Shield_PIO_B_gpio_translator:uav_readdatavalid -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Shield_PIO_B_gpio_translator:uav_debugaccess
	wire   [3:0] shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:m0_byteenable -> Shield_PIO_B_gpio_translator:uav_byteenable
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rf_source_valid -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_data;             // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rf_source_data -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sam9_m1_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // SAM9_M1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         sam9_m1_translator_avalon_universal_master_0_agent_cp_valid;                            // SAM9_M1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         sam9_m1_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // SAM9_M1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [86:0] sam9_m1_translator_avalon_universal_master_0_agent_cp_data;                             // SAM9_M1_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         sam9_m1_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router:sink_ready -> SAM9_M1_translator_avalon_universal_master_0_agent:cp_ready
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_valid;                         // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [86:0] sysid_sysid_translator_avalon_universal_slave_0_agent_rp_data;                          // SysID_SysID_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         sysid_sysid_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router:sink_ready -> SysID_SysID_translator_avalon_universal_slave_0_agent:rp_ready
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                      // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [86:0] funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_data;                       // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_001:sink_ready -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                      // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [86:0] funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_data;                       // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_002:sink_ready -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                      // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [86:0] funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_data;                       // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_003:sink_ready -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                      // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [86:0] funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_data;                       // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_004:sink_ready -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [86:0] shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_005:sink_ready -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [86:0] shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_data;                    // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_006:sink_ready -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:rp_ready
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_valid;                   // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [86:0] shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_data;                    // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_007:sink_ready -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                            // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                  // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                          // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [86:0] addr_router_src_data;                                                                   // addr_router:src_data -> limiter:cmd_sink_data
	wire   [7:0] addr_router_src_channel;                                                                // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                  // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                            // limiter:rsp_src_endofpacket -> SAM9_M1_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                  // limiter:rsp_src_valid -> SAM9_M1_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                          // limiter:rsp_src_startofpacket -> SAM9_M1_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [86:0] limiter_rsp_src_data;                                                                   // limiter:rsp_src_data -> SAM9_M1_translator_avalon_universal_master_0_agent:rp_data
	wire   [7:0] limiter_rsp_src_channel;                                                                // limiter:rsp_src_channel -> SAM9_M1_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                  // SAM9_M1_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         cmd_xbar_demux_src0_endofpacket;                                                        // cmd_xbar_demux:src0_endofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                              // cmd_xbar_demux:src0_valid -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                      // cmd_xbar_demux:src0_startofpacket -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src0_data;                                                               // cmd_xbar_demux:src0_data -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_data
	wire   [7:0] cmd_xbar_demux_src0_channel;                                                            // cmd_xbar_demux:src0_channel -> SysID_SysID_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src1_endofpacket;                                                        // cmd_xbar_demux:src1_endofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                              // cmd_xbar_demux:src1_valid -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                      // cmd_xbar_demux:src1_startofpacket -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src1_data;                                                               // cmd_xbar_demux:src1_data -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire   [7:0] cmd_xbar_demux_src1_channel;                                                            // cmd_xbar_demux:src1_channel -> FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src2_endofpacket;                                                        // cmd_xbar_demux:src2_endofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                              // cmd_xbar_demux:src2_valid -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                      // cmd_xbar_demux:src2_startofpacket -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src2_data;                                                               // cmd_xbar_demux:src2_data -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire   [7:0] cmd_xbar_demux_src2_channel;                                                            // cmd_xbar_demux:src2_channel -> FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src3_endofpacket;                                                        // cmd_xbar_demux:src3_endofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                              // cmd_xbar_demux:src3_valid -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                      // cmd_xbar_demux:src3_startofpacket -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src3_data;                                                               // cmd_xbar_demux:src3_data -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire   [7:0] cmd_xbar_demux_src3_channel;                                                            // cmd_xbar_demux:src3_channel -> FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src4_endofpacket;                                                        // cmd_xbar_demux:src4_endofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                              // cmd_xbar_demux:src4_valid -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                      // cmd_xbar_demux:src4_startofpacket -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src4_data;                                                               // cmd_xbar_demux:src4_data -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire   [7:0] cmd_xbar_demux_src4_channel;                                                            // cmd_xbar_demux:src4_channel -> FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src5_endofpacket;                                                        // cmd_xbar_demux:src5_endofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src5_valid;                                                              // cmd_xbar_demux:src5_valid -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src5_startofpacket;                                                      // cmd_xbar_demux:src5_startofpacket -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src5_data;                                                               // cmd_xbar_demux:src5_data -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire   [7:0] cmd_xbar_demux_src5_channel;                                                            // cmd_xbar_demux:src5_channel -> Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src6_endofpacket;                                                        // cmd_xbar_demux:src6_endofpacket -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src6_valid;                                                              // cmd_xbar_demux:src6_valid -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src6_startofpacket;                                                      // cmd_xbar_demux:src6_startofpacket -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src6_data;                                                               // cmd_xbar_demux:src6_data -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:cp_data
	wire   [7:0] cmd_xbar_demux_src6_channel;                                                            // cmd_xbar_demux:src6_channel -> Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src7_endofpacket;                                                        // cmd_xbar_demux:src7_endofpacket -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src7_valid;                                                              // cmd_xbar_demux:src7_valid -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src7_startofpacket;                                                      // cmd_xbar_demux:src7_startofpacket -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src7_data;                                                               // cmd_xbar_demux:src7_data -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:cp_data
	wire   [7:0] cmd_xbar_demux_src7_channel;                                                            // cmd_xbar_demux:src7_channel -> Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                        // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                              // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                      // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [86:0] rsp_xbar_demux_src0_data;                                                               // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [7:0] rsp_xbar_demux_src0_channel;                                                            // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                              // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                    // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                          // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                  // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [86:0] rsp_xbar_demux_001_src0_data;                                                           // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [7:0] rsp_xbar_demux_001_src0_channel;                                                        // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                          // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                    // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                          // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                  // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [86:0] rsp_xbar_demux_002_src0_data;                                                           // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [7:0] rsp_xbar_demux_002_src0_channel;                                                        // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                          // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                    // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                          // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                  // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [86:0] rsp_xbar_demux_003_src0_data;                                                           // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [7:0] rsp_xbar_demux_003_src0_channel;                                                        // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                          // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                    // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                          // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                  // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [86:0] rsp_xbar_demux_004_src0_data;                                                           // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [7:0] rsp_xbar_demux_004_src0_channel;                                                        // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                          // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                    // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                          // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                  // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [86:0] rsp_xbar_demux_005_src0_data;                                                           // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [7:0] rsp_xbar_demux_005_src0_channel;                                                        // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                          // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                    // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                          // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                  // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [86:0] rsp_xbar_demux_006_src0_data;                                                           // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire   [7:0] rsp_xbar_demux_006_src0_channel;                                                        // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                          // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                    // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                          // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                  // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire  [86:0] rsp_xbar_demux_007_src0_data;                                                           // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire   [7:0] rsp_xbar_demux_007_src0_channel;                                                        // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                          // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                            // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                          // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [86:0] limiter_cmd_src_data;                                                                   // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [7:0] limiter_cmd_src_channel;                                                                // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                  // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                           // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                 // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                         // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [86:0] rsp_xbar_mux_src_data;                                                                  // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [7:0] rsp_xbar_mux_src_channel;                                                               // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                 // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         cmd_xbar_demux_src0_ready;                                                              // SysID_SysID_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire         id_router_src_endofpacket;                                                              // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                    // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                            // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [86:0] id_router_src_data;                                                                     // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [7:0] id_router_src_channel;                                                                  // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                    // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_demux_src1_ready;                                                              // FuncLED_0_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire         id_router_001_src_endofpacket;                                                          // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                        // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [86:0] id_router_001_src_data;                                                                 // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [7:0] id_router_001_src_channel;                                                              // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_src2_ready;                                                              // FuncLED_1_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	wire         id_router_002_src_endofpacket;                                                          // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                        // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [86:0] id_router_002_src_data;                                                                 // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [7:0] id_router_002_src_channel;                                                              // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_src3_ready;                                                              // FuncLED_2_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src3_ready
	wire         id_router_003_src_endofpacket;                                                          // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                        // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [86:0] id_router_003_src_data;                                                                 // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [7:0] id_router_003_src_channel;                                                              // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_src4_ready;                                                              // FuncLED_3_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src4_ready
	wire         id_router_004_src_endofpacket;                                                          // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                        // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [86:0] id_router_004_src_data;                                                                 // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [7:0] id_router_004_src_channel;                                                              // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_src5_ready;                                                              // Shield_Admin_Ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src5_ready
	wire         id_router_005_src_endofpacket;                                                          // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                        // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [86:0] id_router_005_src_data;                                                                 // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [7:0] id_router_005_src_channel;                                                              // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_src6_ready;                                                              // Shield_PIO_A_gpio_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src6_ready
	wire         id_router_006_src_endofpacket;                                                          // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                        // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [86:0] id_router_006_src_data;                                                                 // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [7:0] id_router_006_src_channel;                                                              // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_src7_ready;                                                              // Shield_PIO_B_gpio_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src7_ready
	wire         id_router_007_src_endofpacket;                                                          // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                        // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [86:0] id_router_007_src_data;                                                                 // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [7:0] id_router_007_src_channel;                                                              // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire   [7:0] limiter_cmd_valid_data;                                                                 // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire         irq_mapper_receiver0_irq;                                                               // Shield_Admin:ins_OC_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                               // Shield_PIO_A:ins_INTRQ_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                               // Shield_PIO_B:ins_INTRQ_irq -> irq_mapper:receiver2_irq
	wire   [9:0] sam9_events_irq;                                                                        // irq_synchronizer:sender_irq -> SAM9:inr_EVENTS_irq
	wire   [9:0] irq_synchronizer_receiver_irq;                                                          // irq_mapper:sender_irq -> irq_synchronizer:receiver_irq

	qsys_tabby_host sam9 (
		.rso_MRST_reset       (sam9_mrst_reset),       //   MRST.reset
		.cso_MCLK_clk         (sam9_mclk_clk),         //   MCLK.clk
		.cso_H1CLK_clk        (),                      //  H1CLK.clk
		.cso_H2CLK_clk        (),                      //  H2CLK.clk
		.avm_M1_writedata     (sam9_m1_writedata),     //     M1.writedata
		.avm_M1_readdata      (sam9_m1_readdata),      //       .readdata
		.avm_M1_address       (sam9_m1_address),       //       .address
		.avm_M1_byteenable    (sam9_m1_byteenable),    //       .byteenable
		.avm_M1_write         (sam9_m1_write),         //       .write
		.avm_M1_read          (sam9_m1_read),          //       .read
		.avm_M1_begintransfer (sam9_m1_begintransfer), //       .begintransfer
		.avm_M1_readdatavalid (sam9_m1_readdatavalid), //       .readdatavalid
		.avm_M1_waitrequest   (sam9_m1_waitrequest),   //       .waitrequest
		.inr_EVENTS_irq       (sam9_events_irq),       // EVENTS.irq
		.coe_M1_RSTN          (m1_RSTN),               // EXPORT.export
		.coe_M1_CLK           (m1_CLK),                //       .export
		.coe_M1_ADDR          (m1_ADDR),               //       .export
		.coe_M1_DATA          (m1_DATA),               //       .export
		.coe_M1_CSN           (m1_CSN),                //       .export
		.coe_M1_BEN           (m1_BEN),                //       .export
		.coe_M1_RDN           (m1_RDN),                //       .export
		.coe_M1_WRN           (m1_WRN),                //       .export
		.coe_M1_WAITN         (m1_WAITN),              //       .export
		.coe_M1_EINT          (m1_EINT)                //       .export
	);

	qsys_basic_SysID sysid (
		.rsi_MRST_reset        (sam9_mrst_reset),                                        //  MRST.reset
		.csi_MCLK_clk          (sam9_mclk_clk),                                          //  MCLK.clk
		.avs_SysID_readdata    (sysid_sysid_translator_avalon_anti_slave_0_readdata),    // SysID.readdata
		.avs_SysID_read        (sysid_sysid_translator_avalon_anti_slave_0_read),        //      .read
		.avs_SysID_waitrequest (sysid_sysid_translator_avalon_anti_slave_0_waitrequest)  //      .waitrequest
	);

	qsys_basic_FuncLED funcled_0 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                           //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                             //   MCLK.clk
		.avs_LEDD_writedata   (funcled_0_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (funcled_0_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (funcled_0_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (funcled_0_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (funcled_0_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (funcled_0_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (test_ledstate_0_leds_data),                                 //   LEDS.data
		.asi_LEDS_valid       (test_ledstate_0_leds_valid),                                //       .valid
		.asi_LEDS_ready       (test_ledstate_0_leds_ready),                                //       .ready
		.coe_LED_R            (led_f0_R),                                                  // EXPORT.export
		.coe_LED_G            (led_f0_G),                                                  //       .export
		.coe_LED_B            (led_f0_B)                                                   //       .export
	);

	qsys_basic_FuncLED funcled_1 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                           //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                             //   MCLK.clk
		.avs_LEDD_writedata   (funcled_1_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (funcled_1_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (funcled_1_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (funcled_1_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (funcled_1_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (funcled_1_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (test_ledstate_1_leds_data),                                 //   LEDS.data
		.asi_LEDS_valid       (test_ledstate_1_leds_valid),                                //       .valid
		.asi_LEDS_ready       (test_ledstate_1_leds_ready),                                //       .ready
		.coe_LED_R            (led_f1_R),                                                  // EXPORT.export
		.coe_LED_G            (led_f1_G),                                                  //       .export
		.coe_LED_B            (led_f1_B)                                                   //       .export
	);

	qsys_basic_FuncLED funcled_2 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                           //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                             //   MCLK.clk
		.avs_LEDD_writedata   (funcled_2_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (funcled_2_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (funcled_2_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (funcled_2_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (funcled_2_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (funcled_2_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (test_ledstate_2_leds_data),                                 //   LEDS.data
		.asi_LEDS_valid       (test_ledstate_2_leds_valid),                                //       .valid
		.asi_LEDS_ready       (test_ledstate_2_leds_ready),                                //       .ready
		.coe_LED_R            (led_f2_R),                                                  // EXPORT.export
		.coe_LED_G            (led_f2_G),                                                  //       .export
		.coe_LED_B            (led_f2_B)                                                   //       .export
	);

	qsys_basic_FuncLED funcled_3 (
		.rsi_MRST_reset       (sam9_mrst_reset),                                           //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                             //   MCLK.clk
		.avs_LEDD_writedata   (funcled_3_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (funcled_3_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (funcled_3_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (funcled_3_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (funcled_3_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (funcled_3_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (test_ledstate_3_leds_data),                                 //   LEDS.data
		.asi_LEDS_valid       (test_ledstate_3_leds_valid),                                //       .valid
		.asi_LEDS_ready       (test_ledstate_3_leds_ready),                                //       .ready
		.coe_LED_R            (led_f3_R),                                                  // EXPORT.export
		.coe_LED_G            (led_f3_G),                                                  //       .export
		.coe_LED_B            (led_f3_B)                                                   //       .export
	);

	qsys_shield_moduleBasicCtrl shield_admin (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_Ctrl_writedata   (shield_admin_ctrl_translator_avalon_anti_slave_0_writedata),   //   Ctrl.writedata
		.avs_Ctrl_readdata    (shield_admin_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_Ctrl_byteenable  (shield_admin_ctrl_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_Ctrl_write       (shield_admin_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_Ctrl_read        (shield_admin_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_Ctrl_waitrequest (shield_admin_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.ins_OC_irq           (irq_mapper_receiver0_irq),                                     //     OC.irq
		.coe_A_OCN            (shield_A_OCN),                                                 // EXPORT.export
		.coe_A_PWREN          (shield_A_PWREN),                                               //       .export
		.coe_A_HOE            (shield_A_HOE),                                                 //       .export
		.coe_A_LOE            (shield_A_LOE),                                                 //       .export
		.coe_B_OCN            (shield_B_OCN),                                                 //       .export
		.coe_B_PWREN          (shield_B_PWREN),                                               //       .export
		.coe_B_HOE            (shield_B_HOE),                                                 //       .export
		.coe_B_LOE            (shield_B_LOE)                                                  //       .export
	);

	qsys_test_LEDState test_ledstate_1 (
		.rsi_MRST_reset (sam9_mrst_reset),            // MRST.reset
		.csi_MCLK_clk   (sam9_mclk_clk),              // MCLK.clk
		.aso_LEDS_data  (test_ledstate_1_leds_data),  // LEDS.data
		.aso_LEDS_valid (test_ledstate_1_leds_valid), //     .valid
		.aso_LEDS_ready (test_ledstate_1_leds_ready)  //     .ready
	);

	qsys_test_LEDState test_ledstate_2 (
		.rsi_MRST_reset (sam9_mrst_reset),            // MRST.reset
		.csi_MCLK_clk   (sam9_mclk_clk),              // MCLK.clk
		.aso_LEDS_data  (test_ledstate_2_leds_data),  // LEDS.data
		.aso_LEDS_valid (test_ledstate_2_leds_valid), //     .valid
		.aso_LEDS_ready (test_ledstate_2_leds_ready)  //     .ready
	);

	qsys_test_LEDState test_ledstate_3 (
		.rsi_MRST_reset (sam9_mrst_reset),            // MRST.reset
		.csi_MCLK_clk   (sam9_mclk_clk),              // MCLK.clk
		.aso_LEDS_data  (test_ledstate_3_leds_data),  // LEDS.data
		.aso_LEDS_valid (test_ledstate_3_leds_valid), //     .valid
		.aso_LEDS_ready (test_ledstate_3_leds_ready)  //     .ready
	);

	qsys_test_LEDState test_ledstate_0 (
		.rsi_MRST_reset (sam9_mrst_reset),            // MRST.reset
		.csi_MCLK_clk   (sam9_mclk_clk),              // MCLK.clk
		.aso_LEDS_data  (test_ledstate_0_leds_data),  // LEDS.data
		.aso_LEDS_valid (test_ledstate_0_leds_valid), //     .valid
		.aso_LEDS_ready (test_ledstate_0_leds_ready)  //     .ready
	);

	qsys_shield_pio26b shield_pio_a (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_gpio_writedata   (shield_pio_a_gpio_translator_avalon_anti_slave_0_writedata),   //   gpio.writedata
		.avs_gpio_readdata    (shield_pio_a_gpio_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_gpio_address     (shield_pio_a_gpio_translator_avalon_anti_slave_0_address),     //       .address
		.avs_gpio_byteenable  (shield_pio_a_gpio_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_gpio_write       (shield_pio_a_gpio_translator_avalon_anti_slave_0_write),       //       .write
		.avs_gpio_read        (shield_pio_a_gpio_translator_avalon_anti_slave_0_read),        //       .read
		.avs_gpio_waitrequest (shield_pio_a_gpio_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.ins_INTRQ_irq        (irq_mapper_receiver1_irq),                                     //  INTRQ.irq
		.coe_P0               (slot_a_P0),                                                    // EXPORT.export
		.coe_P1               (slot_a_P1),                                                    //       .export
		.coe_P2               (slot_a_P2),                                                    //       .export
		.coe_P3               (slot_a_P3),                                                    //       .export
		.coe_P4               (slot_a_P4),                                                    //       .export
		.coe_P5               (slot_a_P5),                                                    //       .export
		.coe_P6               (slot_a_P6),                                                    //       .export
		.coe_P7               (slot_a_P7),                                                    //       .export
		.coe_P8               (slot_a_P8),                                                    //       .export
		.coe_P9               (slot_a_P9),                                                    //       .export
		.coe_P10              (slot_a_P10),                                                   //       .export
		.coe_P11              (slot_a_P11),                                                   //       .export
		.coe_P12              (slot_a_P12),                                                   //       .export
		.coe_P13              (slot_a_P13),                                                   //       .export
		.coe_P14              (slot_a_P14),                                                   //       .export
		.coe_P15              (slot_a_P15),                                                   //       .export
		.coe_P16              (slot_a_P16),                                                   //       .export
		.coe_P17              (slot_a_P17),                                                   //       .export
		.coe_P18              (slot_a_P18),                                                   //       .export
		.coe_P19              (slot_a_P19),                                                   //       .export
		.coe_P20              (slot_a_P20),                                                   //       .export
		.coe_P21              (slot_a_P21),                                                   //       .export
		.coe_P22              (slot_a_P22),                                                   //       .export
		.coe_P23              (slot_a_P23),                                                   //       .export
		.coe_P24              (slot_a_P24),                                                   //       .export
		.coe_P25              (slot_a_P25)                                                    //       .export
	);

	qsys_shield_pio26b shield_pio_b (
		.rsi_MRST_reset       (sam9_mrst_reset),                                              //   MRST.reset
		.csi_MCLK_clk         (sam9_mclk_clk),                                                //   MCLK.clk
		.avs_gpio_writedata   (shield_pio_b_gpio_translator_avalon_anti_slave_0_writedata),   //   gpio.writedata
		.avs_gpio_readdata    (shield_pio_b_gpio_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_gpio_address     (shield_pio_b_gpio_translator_avalon_anti_slave_0_address),     //       .address
		.avs_gpio_byteenable  (shield_pio_b_gpio_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_gpio_write       (shield_pio_b_gpio_translator_avalon_anti_slave_0_write),       //       .write
		.avs_gpio_read        (shield_pio_b_gpio_translator_avalon_anti_slave_0_read),        //       .read
		.avs_gpio_waitrequest (shield_pio_b_gpio_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.ins_INTRQ_irq        (irq_mapper_receiver2_irq),                                     //  INTRQ.irq
		.coe_P0               (slot_b_P0),                                                    // EXPORT.export
		.coe_P1               (slot_b_P1),                                                    //       .export
		.coe_P2               (slot_b_P2),                                                    //       .export
		.coe_P3               (slot_b_P3),                                                    //       .export
		.coe_P4               (slot_b_P4),                                                    //       .export
		.coe_P5               (slot_b_P5),                                                    //       .export
		.coe_P6               (slot_b_P6),                                                    //       .export
		.coe_P7               (slot_b_P7),                                                    //       .export
		.coe_P8               (slot_b_P8),                                                    //       .export
		.coe_P9               (slot_b_P9),                                                    //       .export
		.coe_P10              (slot_b_P10),                                                   //       .export
		.coe_P11              (slot_b_P11),                                                   //       .export
		.coe_P12              (slot_b_P12),                                                   //       .export
		.coe_P13              (slot_b_P13),                                                   //       .export
		.coe_P14              (slot_b_P14),                                                   //       .export
		.coe_P15              (slot_b_P15),                                                   //       .export
		.coe_P16              (slot_b_P16),                                                   //       .export
		.coe_P17              (slot_b_P17),                                                   //       .export
		.coe_P18              (slot_b_P18),                                                   //       .export
		.coe_P19              (slot_b_P19),                                                   //       .export
		.coe_P20              (slot_b_P20),                                                   //       .export
		.coe_P21              (slot_b_P21),                                                   //       .export
		.coe_P22              (slot_b_P22),                                                   //       .export
		.coe_P23              (slot_b_P23),                                                   //       .export
		.coe_P24              (slot_b_P24),                                                   //       .export
		.coe_P25              (slot_b_P25)                                                    //       .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (1),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sam9_m1_translator (
		.clk                   (sam9_mclk_clk),                                              //                       clk.clk
		.reset                 (sam9_mrst_reset),                                            //                     reset.reset
		.uav_address           (sam9_m1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sam9_m1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sam9_m1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sam9_m1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sam9_m1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sam9_m1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sam9_m1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sam9_m1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sam9_m1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sam9_m1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sam9_m1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sam9_m1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sam9_m1_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (sam9_m1_byteenable),                                         //                          .byteenable
		.av_begintransfer      (sam9_m1_begintransfer),                                      //                          .begintransfer
		.av_read               (sam9_m1_read),                                               //                          .read
		.av_readdata           (sam9_m1_readdata),                                           //                          .readdata
		.av_readdatavalid      (sam9_m1_readdatavalid),                                      //                          .readdatavalid
		.av_write              (sam9_m1_write),                                              //                          .write
		.av_writedata          (sam9_m1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                       //               (terminated)
		.av_beginbursttransfer (1'b0),                                                       //               (terminated)
		.av_chipselect         (1'b0),                                                       //               (terminated)
		.av_lock               (1'b0),                                                       //               (terminated)
		.av_debugaccess        (1'b0),                                                       //               (terminated)
		.uav_clken             (),                                                           //               (terminated)
		.av_clken              (1'b1)                                                        //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_sysid_translator (
		.clk                   (sam9_mclk_clk),                                                          //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                        //                    reset.reset
		.uav_address           (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read               (sysid_sysid_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata           (sysid_sysid_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_waitrequest        (sysid_sysid_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                       //              (terminated)
		.av_write              (),                                                                       //              (terminated)
		.av_writedata          (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_chipselect         (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) funcled_0_ledd_translator (
		.clk                   (sam9_mclk_clk),                                                             //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                           //                    reset.reset
		.uav_address           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (funcled_0_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (funcled_0_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (funcled_0_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (funcled_0_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (funcled_0_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (funcled_0_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_chipselect         (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) funcled_1_ledd_translator (
		.clk                   (sam9_mclk_clk),                                                             //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                           //                    reset.reset
		.uav_address           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (funcled_1_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (funcled_1_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (funcled_1_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (funcled_1_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (funcled_1_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (funcled_1_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_chipselect         (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) funcled_2_ledd_translator (
		.clk                   (sam9_mclk_clk),                                                             //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                           //                    reset.reset
		.uav_address           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (funcled_2_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (funcled_2_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (funcled_2_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (funcled_2_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (funcled_2_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (funcled_2_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_chipselect         (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) funcled_3_ledd_translator (
		.clk                   (sam9_mclk_clk),                                                             //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                           //                    reset.reset
		.uav_address           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (funcled_3_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (funcled_3_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (funcled_3_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (funcled_3_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (funcled_3_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (funcled_3_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_chipselect         (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shield_admin_ctrl_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (shield_admin_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (shield_admin_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shield_admin_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shield_admin_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (shield_admin_ctrl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (shield_admin_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shield_pio_a_gpio_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (shield_pio_a_gpio_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (shield_pio_a_gpio_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (shield_pio_a_gpio_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shield_pio_a_gpio_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shield_pio_a_gpio_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (shield_pio_a_gpio_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (shield_pio_a_gpio_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) shield_pio_b_gpio_translator (
		.clk                   (sam9_mclk_clk),                                                                //                      clk.clk
		.reset                 (sam9_mrst_reset),                                                              //                    reset.reset
		.uav_address           (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (shield_pio_b_gpio_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (shield_pio_b_gpio_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (shield_pio_b_gpio_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (shield_pio_b_gpio_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (shield_pio_b_gpio_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (shield_pio_b_gpio_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (shield_pio_b_gpio_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) funcled_0_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                       //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                     //       clk_reset.reset
		.m0_address              (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (funcled_0_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                         //                .channel
		.rf_sink_ready           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                       //       clk.clk
		.reset             (sam9_mrst_reset),                                                                     // clk_reset.reset
		.in_data           (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_sysid_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                    //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                  //       clk_reset.reset
		.m0_address              (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_sysid_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                      //                .channel
		.rf_sink_ready           (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_sysid_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                    //       clk.clk
		.reset             (sam9_mrst_reset),                                                                  // clk_reset.reset
		.in_data           (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_sysid_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (8),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7)
	) sam9_m1_translator_avalon_universal_master_0_agent (
		.clk              (sam9_mclk_clk),                                                       //       clk.clk
		.reset            (sam9_mrst_reset),                                                     // clk_reset.reset
		.av_address       (sam9_m1_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sam9_m1_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sam9_m1_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sam9_m1_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sam9_m1_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sam9_m1_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sam9_m1_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sam9_m1_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sam9_m1_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sam9_m1_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sam9_m1_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sam9_m1_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sam9_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sam9_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sam9_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sam9_m1_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                               //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                //          .data
		.rp_channel       (limiter_rsp_src_channel),                                             //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                       //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                         //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shield_pio_a_gpio_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src6_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_src6_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_src6_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_src6_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src6_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src6_channel),                                                            //                .channel
		.rf_sink_ready           (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) funcled_3_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                       //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                     //       clk_reset.reset
		.m0_address              (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (funcled_3_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src4_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_src4_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_src4_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_src4_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src4_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src4_channel),                                                         //                .channel
		.rf_sink_ready           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                       //       clk.clk
		.reset             (sam9_mrst_reset),                                                                     // clk_reset.reset
		.in_data           (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shield_admin_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src5_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_src5_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_src5_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_src5_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src5_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src5_channel),                                                            //                .channel
		.rf_sink_ready           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) funcled_2_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                       //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                     //       clk_reset.reset
		.m0_address              (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (funcled_2_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src3_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_src3_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_src3_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_src3_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src3_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src3_channel),                                                         //                .channel
		.rf_sink_ready           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                       //       clk.clk
		.reset             (sam9_mrst_reset),                                                                     // clk_reset.reset
		.in_data           (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) funcled_1_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                       //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                     //       clk_reset.reset
		.m0_address              (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (funcled_1_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src2_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_src2_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_src2_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_src2_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src2_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src2_channel),                                                         //                .channel
		.rf_sink_ready           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                       //       clk.clk
		.reset             (sam9_mrst_reset),                                                                     // clk_reset.reset
		.in_data           (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) shield_pio_b_gpio_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_mclk_clk),                                                                          //             clk.clk
		.reset                   (sam9_mrst_reset),                                                                        //       clk_reset.reset
		.m0_address              (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src7_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_src7_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_src7_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_src7_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src7_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src7_channel),                                                            //                .channel
		.rf_sink_ready           (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_mclk_clk),                                                                          //       clk.clk
		.reset             (sam9_mrst_reset),                                                                        // clk_reset.reset
		.in_data           (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	frontier_addr_router addr_router (
		.sink_ready         (sam9_m1_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sam9_m1_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sam9_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sam9_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sam9_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                       //       clk.clk
		.reset              (sam9_mrst_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                               //       src.ready
		.src_valid          (addr_router_src_valid),                                               //          .valid
		.src_data           (addr_router_src_data),                                                //          .data
		.src_channel        (addr_router_src_channel),                                             //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                          //          .endofpacket
	);

	frontier_id_router id_router (
		.sink_ready         (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_sysid_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                          //       clk.clk
		.reset              (sam9_mrst_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                    //       src.ready
		.src_valid          (id_router_src_valid),                                                    //          .valid
		.src_data           (id_router_src_data),                                                     //          .data
		.src_channel        (id_router_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                               //          .endofpacket
	);

	frontier_id_router id_router_001 (
		.sink_ready         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (funcled_0_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                             //       clk.clk
		.reset              (sam9_mrst_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                   //       src.ready
		.src_valid          (id_router_001_src_valid),                                                   //          .valid
		.src_data           (id_router_001_src_data),                                                    //          .data
		.src_channel        (id_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                              //          .endofpacket
	);

	frontier_id_router id_router_002 (
		.sink_ready         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (funcled_1_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                             //       clk.clk
		.reset              (sam9_mrst_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                   //       src.ready
		.src_valid          (id_router_002_src_valid),                                                   //          .valid
		.src_data           (id_router_002_src_data),                                                    //          .data
		.src_channel        (id_router_002_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                              //          .endofpacket
	);

	frontier_id_router id_router_003 (
		.sink_ready         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (funcled_2_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                             //       clk.clk
		.reset              (sam9_mrst_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                   //       src.ready
		.src_valid          (id_router_003_src_valid),                                                   //          .valid
		.src_data           (id_router_003_src_data),                                                    //          .data
		.src_channel        (id_router_003_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                              //          .endofpacket
	);

	frontier_id_router id_router_004 (
		.sink_ready         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (funcled_3_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                             //       clk.clk
		.reset              (sam9_mrst_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                   //       src.ready
		.src_valid          (id_router_004_src_valid),                                                   //          .valid
		.src_data           (id_router_004_src_data),                                                    //          .data
		.src_channel        (id_router_004_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                              //          .endofpacket
	);

	frontier_id_router id_router_005 (
		.sink_ready         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shield_admin_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                      //       src.ready
		.src_valid          (id_router_005_src_valid),                                                      //          .valid
		.src_data           (id_router_005_src_data),                                                       //          .data
		.src_channel        (id_router_005_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router id_router_006 (
		.sink_ready         (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shield_pio_a_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                      //       src.ready
		.src_valid          (id_router_006_src_valid),                                                      //          .valid
		.src_data           (id_router_006_src_data),                                                       //          .data
		.src_channel        (id_router_006_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router id_router_007 (
		.sink_ready         (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (shield_pio_b_gpio_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_mclk_clk),                                                                //       clk.clk
		.reset              (sam9_mrst_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                      //       src.ready
		.src_valid          (id_router_007_src_valid),                                                      //          .valid
		.src_data           (id_router_007_src_data),                                                       //          .data
		.src_channel        (id_router_007_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                 //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (8),
		.VALID_WIDTH               (8),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (sam9_mclk_clk),                  //       clk.clk
		.reset                  (sam9_mrst_reset),                // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	frontier_cmd_xbar_demux cmd_xbar_demux (
		.clk                (sam9_mclk_clk),                     //        clk.clk
		.reset              (sam9_mrst_reset),                   //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_src6_endofpacket),   //           .endofpacket
		.src7_ready         (cmd_xbar_demux_src7_ready),         //       src7.ready
		.src7_valid         (cmd_xbar_demux_src7_valid),         //           .valid
		.src7_data          (cmd_xbar_demux_src7_data),          //           .data
		.src7_channel       (cmd_xbar_demux_src7_channel),       //           .channel
		.src7_startofpacket (cmd_xbar_demux_src7_startofpacket), //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_src7_endofpacket)    //           .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux (
		.clk                (sam9_mclk_clk),                     //       clk.clk
		.reset              (sam9_mrst_reset),                   // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_007 (
		.clk                (sam9_mclk_clk),                         //       clk.clk
		.reset              (sam9_mrst_reset),                       // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (sam9_mclk_clk),                         //       clk.clk
		.reset               (sam9_mrst_reset),                       // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	frontier_irq_mapper irq_mapper (
		.clk           (sam9_mclk_clk),                 //       clk.clk
		.reset         (sam9_mrst_reset),               // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),      // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),      // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),      // receiver2.irq
		.sender_irq    (irq_synchronizer_receiver_irq)  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (10)
	) irq_synchronizer (
		.receiver_clk   (sam9_mclk_clk),                 //       receiver_clk.clk
		.sender_clk     (sam9_mclk_clk),                 //         sender_clk.clk
		.receiver_reset (sam9_mrst_reset),               // receiver_clk_reset.reset
		.sender_reset   (sam9_mrst_reset),               //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq), //           receiver.irq
		.sender_irq     (sam9_events_irq)                //             sender.irq
	);

endmodule
