// frontier.v

// Generated using ACDS version 11.1sp2 259 at 2012.07.18.19:01:15

`timescale 1 ps / 1 ps
module frontier (
		output wire        led_f3_R,      // led_f3.R
		output wire        led_f3_G,      //       .G
		output wire        led_f3_B,      //       .B
		output wire        led_f2_R,      // led_f2.R
		output wire        led_f2_G,      //       .G
		output wire        led_f2_B,      //       .B
		input  wire        admin_A_OCN,   //  admin.A_OCN
		output wire        admin_A_PWREN, //       .A_PWREN
		output wire        admin_A_HOE,   //       .A_HOE
		output wire        admin_A_LOE,   //       .A_LOE
		input  wire        admin_B_OCN,   //       .B_OCN
		output wire        admin_B_PWREN, //       .B_PWREN
		output wire        admin_B_HOE,   //       .B_HOE
		output wire        admin_B_LOE,   //       .B_LOE
		input  wire        m1_RSTN,       //     m1.RSTN
		input  wire        m1_CLK,        //       .CLK
		input  wire [21:0] m1_ADDR,       //       .ADDR
		inout  wire [31:0] m1_DATA,       //       .DATA
		input  wire [3:0]  m1_CSN,        //       .CSN
		input  wire [3:0]  m1_BEN,        //       .BEN
		input  wire        m1_RDN,        //       .RDN
		input  wire        m1_WRN,        //       .WRN
		output wire        m1_WAITN,      //       .WAITN
		output wire [9:0]  m1_EINT,       //       .EINT
		output wire        led_f0_R,      // led_f0.R
		output wire        led_f0_G,      //       .G
		output wire        led_f0_B,      //       .B
		output wire        led_f1_R,      // led_f1.R
		output wire        led_f1_G,      //       .G
		output wire        led_f1_B       //       .B
	);

	wire         sam9_host_mrst_reset;                                                                                       // SAM9_HOST:rso_MRST_reset -> [RGB_LED_F0:rsi_MRST_reset, RGB_LED_F0S:rsi_MRST_reset, RGB_LED_F0_LEDD_translator:reset, RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:reset, RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RGB_LED_F1:rsi_MRST_reset, RGB_LED_F1S:rsi_MRST_reset, RGB_LED_F1_LEDD_translator:reset, RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:reset, RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RGB_LED_F2:rsi_MRST_reset, RGB_LED_F2S:rsi_MRST_reset, RGB_LED_F2_LEDD_translator:reset, RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:reset, RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RGB_LED_F3:rsi_MRST_reset, RGB_LED_F3S:rsi_MRST_reset, RGB_LED_F3_LEDD_translator:reset, RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:reset, RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SAM9_HOST_M1_translator:reset, SAM9_HOST_M1_translator_avalon_universal_master_0_agent:reset, TEST_REG_0:rsi_MRST_reset, TEST_REG_0_TestReg_translator:reset, TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:reset, TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, cmd_xbar_demux:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, irq_mapper:reset, irq_synchronizer:receiver_reset, irq_synchronizer:sender_reset, limiter:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, qsys_basic_lophilo_module_ctrl_0:rsi_MRST_reset, qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:reset, qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:reset, qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_mux:reset]
	wire         sam9_host_mclk_clk;                                                                                         // SAM9_HOST:cso_MCLK_clk -> [RGB_LED_F0:csi_MCLK_clk, RGB_LED_F0S:csi_MCLK_clk, RGB_LED_F0_LEDD_translator:clk, RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:clk, RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, RGB_LED_F1:csi_MCLK_clk, RGB_LED_F1S:csi_MCLK_clk, RGB_LED_F1_LEDD_translator:clk, RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:clk, RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, RGB_LED_F2:csi_MCLK_clk, RGB_LED_F2S:csi_MCLK_clk, RGB_LED_F2_LEDD_translator:clk, RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:clk, RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, RGB_LED_F3:csi_MCLK_clk, RGB_LED_F3S:csi_MCLK_clk, RGB_LED_F3_LEDD_translator:clk, RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:clk, RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, SAM9_HOST_M1_translator:clk, SAM9_HOST_M1_translator_avalon_universal_master_0_agent:clk, TEST_REG_0:csi_MCLK_clk, TEST_REG_0_TestReg_translator:clk, TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:clk, TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, cmd_xbar_demux:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, irq_mapper:clk, irq_synchronizer:receiver_clk, irq_synchronizer:sender_clk, limiter:clk, onchip_memory2_0:clk, onchip_memory2_0_s1_translator:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, qsys_basic_lophilo_module_ctrl_0:csi_MCLK_clk, qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:clk, qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:clk, qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_mux:clk]
	wire         rgb_led_f0s_leds_valid;                                                                                     // RGB_LED_F0S:aso_LEDS_valid -> RGB_LED_F0:asi_LEDS_valid
	wire  [23:0] rgb_led_f0s_leds_data;                                                                                      // RGB_LED_F0S:aso_LEDS_data -> RGB_LED_F0:asi_LEDS_data
	wire         rgb_led_f0s_leds_ready;                                                                                     // RGB_LED_F0:asi_LEDS_ready -> RGB_LED_F0S:aso_LEDS_ready
	wire         rgb_led_f1s_leds_valid;                                                                                     // RGB_LED_F1S:aso_LEDS_valid -> RGB_LED_F1:asi_LEDS_valid
	wire  [23:0] rgb_led_f1s_leds_data;                                                                                      // RGB_LED_F1S:aso_LEDS_data -> RGB_LED_F1:asi_LEDS_data
	wire         rgb_led_f1s_leds_ready;                                                                                     // RGB_LED_F1:asi_LEDS_ready -> RGB_LED_F1S:aso_LEDS_ready
	wire         rgb_led_f2s_leds_valid;                                                                                     // RGB_LED_F2S:aso_LEDS_valid -> RGB_LED_F2:asi_LEDS_valid
	wire  [23:0] rgb_led_f2s_leds_data;                                                                                      // RGB_LED_F2S:aso_LEDS_data -> RGB_LED_F2:asi_LEDS_data
	wire         rgb_led_f2s_leds_ready;                                                                                     // RGB_LED_F2:asi_LEDS_ready -> RGB_LED_F2S:aso_LEDS_ready
	wire         rgb_led_f3s_leds_valid;                                                                                     // RGB_LED_F3S:aso_LEDS_valid -> RGB_LED_F3:asi_LEDS_valid
	wire  [23:0] rgb_led_f3s_leds_data;                                                                                      // RGB_LED_F3S:aso_LEDS_data -> RGB_LED_F3:asi_LEDS_data
	wire         rgb_led_f3s_leds_ready;                                                                                     // RGB_LED_F3:asi_LEDS_ready -> RGB_LED_F3S:aso_LEDS_ready
	wire         sam9_host_m1_waitrequest;                                                                                   // SAM9_HOST_M1_translator:av_waitrequest -> SAM9_HOST:avm_M1_waitrequest
	wire  [31:0] sam9_host_m1_address;                                                                                       // SAM9_HOST:avm_M1_address -> SAM9_HOST_M1_translator:av_address
	wire  [31:0] sam9_host_m1_writedata;                                                                                     // SAM9_HOST:avm_M1_writedata -> SAM9_HOST_M1_translator:av_writedata
	wire         sam9_host_m1_write;                                                                                         // SAM9_HOST:avm_M1_write -> SAM9_HOST_M1_translator:av_write
	wire         sam9_host_m1_read;                                                                                          // SAM9_HOST:avm_M1_read -> SAM9_HOST_M1_translator:av_read
	wire  [31:0] sam9_host_m1_readdata;                                                                                      // SAM9_HOST_M1_translator:av_readdata -> SAM9_HOST:avm_M1_readdata
	wire         sam9_host_m1_begintransfer;                                                                                 // SAM9_HOST:avm_M1_begintransfer -> SAM9_HOST_M1_translator:av_begintransfer
	wire         sam9_host_m1_readdatavalid;                                                                                 // SAM9_HOST_M1_translator:av_readdatavalid -> SAM9_HOST:avm_M1_readdatavalid
	wire   [3:0] sam9_host_m1_byteenable;                                                                                    // SAM9_HOST:avm_M1_byteenable -> SAM9_HOST_M1_translator:av_byteenable
	wire         rgb_led_f0_ledd_translator_avalon_anti_slave_0_waitrequest;                                                 // RGB_LED_F0:avs_LEDD_waitrequest -> RGB_LED_F0_LEDD_translator:av_waitrequest
	wire  [31:0] rgb_led_f0_ledd_translator_avalon_anti_slave_0_writedata;                                                   // RGB_LED_F0_LEDD_translator:av_writedata -> RGB_LED_F0:avs_LEDD_writedata
	wire         rgb_led_f0_ledd_translator_avalon_anti_slave_0_write;                                                       // RGB_LED_F0_LEDD_translator:av_write -> RGB_LED_F0:avs_LEDD_write
	wire         rgb_led_f0_ledd_translator_avalon_anti_slave_0_read;                                                        // RGB_LED_F0_LEDD_translator:av_read -> RGB_LED_F0:avs_LEDD_read
	wire  [31:0] rgb_led_f0_ledd_translator_avalon_anti_slave_0_readdata;                                                    // RGB_LED_F0:avs_LEDD_readdata -> RGB_LED_F0_LEDD_translator:av_readdata
	wire   [3:0] rgb_led_f0_ledd_translator_avalon_anti_slave_0_byteenable;                                                  // RGB_LED_F0_LEDD_translator:av_byteenable -> RGB_LED_F0:avs_LEDD_byteenable
	wire         rgb_led_f1_ledd_translator_avalon_anti_slave_0_waitrequest;                                                 // RGB_LED_F1:avs_LEDD_waitrequest -> RGB_LED_F1_LEDD_translator:av_waitrequest
	wire  [31:0] rgb_led_f1_ledd_translator_avalon_anti_slave_0_writedata;                                                   // RGB_LED_F1_LEDD_translator:av_writedata -> RGB_LED_F1:avs_LEDD_writedata
	wire         rgb_led_f1_ledd_translator_avalon_anti_slave_0_write;                                                       // RGB_LED_F1_LEDD_translator:av_write -> RGB_LED_F1:avs_LEDD_write
	wire         rgb_led_f1_ledd_translator_avalon_anti_slave_0_read;                                                        // RGB_LED_F1_LEDD_translator:av_read -> RGB_LED_F1:avs_LEDD_read
	wire  [31:0] rgb_led_f1_ledd_translator_avalon_anti_slave_0_readdata;                                                    // RGB_LED_F1:avs_LEDD_readdata -> RGB_LED_F1_LEDD_translator:av_readdata
	wire   [3:0] rgb_led_f1_ledd_translator_avalon_anti_slave_0_byteenable;                                                  // RGB_LED_F1_LEDD_translator:av_byteenable -> RGB_LED_F1:avs_LEDD_byteenable
	wire         rgb_led_f2_ledd_translator_avalon_anti_slave_0_waitrequest;                                                 // RGB_LED_F2:avs_LEDD_waitrequest -> RGB_LED_F2_LEDD_translator:av_waitrequest
	wire  [31:0] rgb_led_f2_ledd_translator_avalon_anti_slave_0_writedata;                                                   // RGB_LED_F2_LEDD_translator:av_writedata -> RGB_LED_F2:avs_LEDD_writedata
	wire         rgb_led_f2_ledd_translator_avalon_anti_slave_0_write;                                                       // RGB_LED_F2_LEDD_translator:av_write -> RGB_LED_F2:avs_LEDD_write
	wire         rgb_led_f2_ledd_translator_avalon_anti_slave_0_read;                                                        // RGB_LED_F2_LEDD_translator:av_read -> RGB_LED_F2:avs_LEDD_read
	wire  [31:0] rgb_led_f2_ledd_translator_avalon_anti_slave_0_readdata;                                                    // RGB_LED_F2:avs_LEDD_readdata -> RGB_LED_F2_LEDD_translator:av_readdata
	wire   [3:0] rgb_led_f2_ledd_translator_avalon_anti_slave_0_byteenable;                                                  // RGB_LED_F2_LEDD_translator:av_byteenable -> RGB_LED_F2:avs_LEDD_byteenable
	wire         rgb_led_f3_ledd_translator_avalon_anti_slave_0_waitrequest;                                                 // RGB_LED_F3:avs_LEDD_waitrequest -> RGB_LED_F3_LEDD_translator:av_waitrequest
	wire  [31:0] rgb_led_f3_ledd_translator_avalon_anti_slave_0_writedata;                                                   // RGB_LED_F3_LEDD_translator:av_writedata -> RGB_LED_F3:avs_LEDD_writedata
	wire         rgb_led_f3_ledd_translator_avalon_anti_slave_0_write;                                                       // RGB_LED_F3_LEDD_translator:av_write -> RGB_LED_F3:avs_LEDD_write
	wire         rgb_led_f3_ledd_translator_avalon_anti_slave_0_read;                                                        // RGB_LED_F3_LEDD_translator:av_read -> RGB_LED_F3:avs_LEDD_read
	wire  [31:0] rgb_led_f3_ledd_translator_avalon_anti_slave_0_readdata;                                                    // RGB_LED_F3:avs_LEDD_readdata -> RGB_LED_F3_LEDD_translator:av_readdata
	wire   [3:0] rgb_led_f3_ledd_translator_avalon_anti_slave_0_byteenable;                                                  // RGB_LED_F3_LEDD_translator:av_byteenable -> RGB_LED_F3:avs_LEDD_byteenable
	wire         test_reg_0_testreg_translator_avalon_anti_slave_0_waitrequest;                                              // TEST_REG_0:avs_TestReg_waitrequest -> TEST_REG_0_TestReg_translator:av_waitrequest
	wire  [31:0] test_reg_0_testreg_translator_avalon_anti_slave_0_writedata;                                                // TEST_REG_0_TestReg_translator:av_writedata -> TEST_REG_0:avs_TestReg_writedata
	wire         test_reg_0_testreg_translator_avalon_anti_slave_0_write;                                                    // TEST_REG_0_TestReg_translator:av_write -> TEST_REG_0:avs_TestReg_write
	wire         test_reg_0_testreg_translator_avalon_anti_slave_0_read;                                                     // TEST_REG_0_TestReg_translator:av_read -> TEST_REG_0:avs_TestReg_read
	wire  [31:0] test_reg_0_testreg_translator_avalon_anti_slave_0_readdata;                                                 // TEST_REG_0:avs_TestReg_readdata -> TEST_REG_0_TestReg_translator:av_readdata
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                               // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire   [9:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                                 // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                              // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                                   // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                                   // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                                // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire   [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                              // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_waitrequest;                           // qsys_basic_lophilo_module_ctrl_0:avs_Ctrl_waitrequest -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:av_waitrequest
	wire  [31:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_writedata;                             // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:av_writedata -> qsys_basic_lophilo_module_ctrl_0:avs_Ctrl_writedata
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_write;                                 // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:av_write -> qsys_basic_lophilo_module_ctrl_0:avs_Ctrl_write
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_read;                                  // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:av_read -> qsys_basic_lophilo_module_ctrl_0:avs_Ctrl_read
	wire  [31:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_readdata;                              // qsys_basic_lophilo_module_ctrl_0:avs_Ctrl_readdata -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:av_readdata
	wire   [3:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_byteenable;                            // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:av_byteenable -> qsys_basic_lophilo_module_ctrl_0:avs_Ctrl_byteenable
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // RGB_LED_F2_LEDD_translator:uav_waitrequest -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> RGB_LED_F2_LEDD_translator:uav_burstcount
	wire  [31:0] rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> RGB_LED_F2_LEDD_translator:uav_writedata
	wire  [31:0] rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_address;                                       // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> RGB_LED_F2_LEDD_translator:uav_address
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_write;                                         // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> RGB_LED_F2_LEDD_translator:uav_write
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                                          // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> RGB_LED_F2_LEDD_translator:uav_lock
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_read;                                          // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> RGB_LED_F2_LEDD_translator:uav_read
	wire  [31:0] rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // RGB_LED_F2_LEDD_translator:uav_readdata -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // RGB_LED_F2_LEDD_translator:uav_readdatavalid -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RGB_LED_F2_LEDD_translator:uav_debugaccess
	wire   [3:0] rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> RGB_LED_F2_LEDD_translator:uav_byteenable
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // RGB_LED_F3_LEDD_translator:uav_waitrequest -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> RGB_LED_F3_LEDD_translator:uav_burstcount
	wire  [31:0] rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> RGB_LED_F3_LEDD_translator:uav_writedata
	wire  [31:0] rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_address;                                       // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> RGB_LED_F3_LEDD_translator:uav_address
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_write;                                         // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> RGB_LED_F3_LEDD_translator:uav_write
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                                          // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> RGB_LED_F3_LEDD_translator:uav_lock
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_read;                                          // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> RGB_LED_F3_LEDD_translator:uav_read
	wire  [31:0] rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // RGB_LED_F3_LEDD_translator:uav_readdata -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // RGB_LED_F3_LEDD_translator:uav_readdatavalid -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RGB_LED_F3_LEDD_translator:uav_debugaccess
	wire   [3:0] rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> RGB_LED_F3_LEDD_translator:uav_byteenable
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // RGB_LED_F0_LEDD_translator:uav_waitrequest -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> RGB_LED_F0_LEDD_translator:uav_burstcount
	wire  [31:0] rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> RGB_LED_F0_LEDD_translator:uav_writedata
	wire  [31:0] rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_address;                                       // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> RGB_LED_F0_LEDD_translator:uav_address
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_write;                                         // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> RGB_LED_F0_LEDD_translator:uav_write
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                                          // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> RGB_LED_F0_LEDD_translator:uav_lock
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_read;                                          // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> RGB_LED_F0_LEDD_translator:uav_read
	wire  [31:0] rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // RGB_LED_F0_LEDD_translator:uav_readdata -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // RGB_LED_F0_LEDD_translator:uav_readdatavalid -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RGB_LED_F0_LEDD_translator:uav_debugaccess
	wire   [3:0] rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> RGB_LED_F0_LEDD_translator:uav_byteenable
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // TEST_REG_0_TestReg_translator:uav_waitrequest -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:m0_burstcount -> TEST_REG_0_TestReg_translator:uav_burstcount
	wire  [31:0] test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:m0_writedata -> TEST_REG_0_TestReg_translator:uav_writedata
	wire  [31:0] test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_address;                                    // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:m0_address -> TEST_REG_0_TestReg_translator:uav_address
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_write;                                      // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:m0_write -> TEST_REG_0_TestReg_translator:uav_write
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_lock;                                       // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:m0_lock -> TEST_REG_0_TestReg_translator:uav_lock
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_read;                                       // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:m0_read -> TEST_REG_0_TestReg_translator:uav_read
	wire  [31:0] test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // TEST_REG_0_TestReg_translator:uav_readdata -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // TEST_REG_0_TestReg_translator:uav_readdatavalid -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:m0_debugaccess -> TEST_REG_0_TestReg_translator:uav_debugaccess
	wire   [3:0] test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:m0_byteenable -> TEST_REG_0_TestReg_translator:uav_byteenable
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rf_source_valid -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_data;                                // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rf_source_data -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_ready -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // RGB_LED_F1_LEDD_translator:uav_waitrequest -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:m0_burstcount -> RGB_LED_F1_LEDD_translator:uav_burstcount
	wire  [31:0] rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:m0_writedata -> RGB_LED_F1_LEDD_translator:uav_writedata
	wire  [31:0] rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_address;                                       // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:m0_address -> RGB_LED_F1_LEDD_translator:uav_address
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_write;                                         // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:m0_write -> RGB_LED_F1_LEDD_translator:uav_write
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_lock;                                          // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:m0_lock -> RGB_LED_F1_LEDD_translator:uav_lock
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_read;                                          // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:m0_read -> RGB_LED_F1_LEDD_translator:uav_read
	wire  [31:0] rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // RGB_LED_F1_LEDD_translator:uav_readdata -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // RGB_LED_F1_LEDD_translator:uav_readdatavalid -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RGB_LED_F1_LEDD_translator:uav_debugaccess
	wire   [3:0] rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:m0_byteenable -> RGB_LED_F1_LEDD_translator:uav_byteenable
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_valid -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_data -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sam9_host_m1_translator_avalon_universal_master_0_waitrequest;                                              // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_waitrequest -> SAM9_HOST_M1_translator:uav_waitrequest
	wire   [2:0] sam9_host_m1_translator_avalon_universal_master_0_burstcount;                                               // SAM9_HOST_M1_translator:uav_burstcount -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] sam9_host_m1_translator_avalon_universal_master_0_writedata;                                                // SAM9_HOST_M1_translator:uav_writedata -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] sam9_host_m1_translator_avalon_universal_master_0_address;                                                  // SAM9_HOST_M1_translator:uav_address -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_address
	wire         sam9_host_m1_translator_avalon_universal_master_0_lock;                                                     // SAM9_HOST_M1_translator:uav_lock -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_lock
	wire         sam9_host_m1_translator_avalon_universal_master_0_write;                                                    // SAM9_HOST_M1_translator:uav_write -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_write
	wire         sam9_host_m1_translator_avalon_universal_master_0_read;                                                     // SAM9_HOST_M1_translator:uav_read -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] sam9_host_m1_translator_avalon_universal_master_0_readdata;                                                 // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_readdata -> SAM9_HOST_M1_translator:uav_readdata
	wire         sam9_host_m1_translator_avalon_universal_master_0_debugaccess;                                              // SAM9_HOST_M1_translator:uav_debugaccess -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] sam9_host_m1_translator_avalon_universal_master_0_byteenable;                                               // SAM9_HOST_M1_translator:uav_byteenable -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_byteenable
	wire         sam9_host_m1_translator_avalon_universal_master_0_readdatavalid;                                            // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_readdatavalid -> SAM9_HOST_M1_translator:uav_readdatavalid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:uav_waitrequest -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:m0_burstcount -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:uav_burstcount
	wire  [31:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata;               // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:m0_writedata -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:uav_writedata
	wire  [31:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address;                 // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:m0_address -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:uav_address
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write;                   // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:m0_write -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:uav_write
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock;                    // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:m0_lock -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:uav_lock
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read;                    // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:m0_read -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:uav_read
	wire  [31:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata;                // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:uav_readdata -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:uav_readdatavalid -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:uav_debugaccess
	wire   [3:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:m0_byteenable -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator:uav_byteenable
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_valid -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data;             // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_data -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sam9_host_m1_translator_avalon_universal_master_0_agent_cp_endofpacket;                                     // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         sam9_host_m1_translator_avalon_universal_master_0_agent_cp_valid;                                           // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         sam9_host_m1_translator_avalon_universal_master_0_agent_cp_startofpacket;                                   // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [86:0] sam9_host_m1_translator_avalon_universal_master_0_agent_cp_data;                                            // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         sam9_host_m1_translator_avalon_universal_master_0_agent_cp_ready;                                           // addr_router:sink_ready -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:cp_ready
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                                         // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [86:0] rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_data;                                          // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router:sink_ready -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                                         // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [86:0] rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_data;                                          // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_001:sink_ready -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                                         // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [86:0] rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_data;                                          // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_002:sink_ready -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_valid;                                         // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [86:0] rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_data;                                          // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_003:sink_ready -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:rp_ready
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_valid;                                      // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [86:0] test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_data;                                       // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_004:sink_ready -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [86:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_005:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid;                   // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [86:0] qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data;                    // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_006:sink_ready -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                                // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                                      // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                              // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [86:0] addr_router_src_data;                                                                                       // addr_router:src_data -> limiter:cmd_sink_data
	wire   [6:0] addr_router_src_channel;                                                                                    // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                                      // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                                // limiter:rsp_src_endofpacket -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                                      // limiter:rsp_src_valid -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                              // limiter:rsp_src_startofpacket -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [86:0] limiter_rsp_src_data;                                                                                       // limiter:rsp_src_data -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_data
	wire   [6:0] limiter_rsp_src_channel;                                                                                    // limiter:rsp_src_channel -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                                      // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         cmd_xbar_demux_src0_endofpacket;                                                                            // cmd_xbar_demux:src0_endofpacket -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                                  // cmd_xbar_demux:src0_valid -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                          // cmd_xbar_demux:src0_startofpacket -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src0_data;                                                                                   // cmd_xbar_demux:src0_data -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src0_channel;                                                                                // cmd_xbar_demux:src0_channel -> RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src1_endofpacket;                                                                            // cmd_xbar_demux:src1_endofpacket -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                                  // cmd_xbar_demux:src1_valid -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                          // cmd_xbar_demux:src1_startofpacket -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src1_data;                                                                                   // cmd_xbar_demux:src1_data -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src1_channel;                                                                                // cmd_xbar_demux:src1_channel -> RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src2_endofpacket;                                                                            // cmd_xbar_demux:src2_endofpacket -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                                  // cmd_xbar_demux:src2_valid -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                          // cmd_xbar_demux:src2_startofpacket -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src2_data;                                                                                   // cmd_xbar_demux:src2_data -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src2_channel;                                                                                // cmd_xbar_demux:src2_channel -> RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src3_endofpacket;                                                                            // cmd_xbar_demux:src3_endofpacket -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                                  // cmd_xbar_demux:src3_valid -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                          // cmd_xbar_demux:src3_startofpacket -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src3_data;                                                                                   // cmd_xbar_demux:src3_data -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src3_channel;                                                                                // cmd_xbar_demux:src3_channel -> RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src4_endofpacket;                                                                            // cmd_xbar_demux:src4_endofpacket -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                                                  // cmd_xbar_demux:src4_valid -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                                          // cmd_xbar_demux:src4_startofpacket -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src4_data;                                                                                   // cmd_xbar_demux:src4_data -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src4_channel;                                                                                // cmd_xbar_demux:src4_channel -> TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src5_endofpacket;                                                                            // cmd_xbar_demux:src5_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src5_valid;                                                                                  // cmd_xbar_demux:src5_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src5_startofpacket;                                                                          // cmd_xbar_demux:src5_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src5_data;                                                                                   // cmd_xbar_demux:src5_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src5_channel;                                                                                // cmd_xbar_demux:src5_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src6_endofpacket;                                                                            // cmd_xbar_demux:src6_endofpacket -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src6_valid;                                                                                  // cmd_xbar_demux:src6_valid -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src6_startofpacket;                                                                          // cmd_xbar_demux:src6_startofpacket -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src6_data;                                                                                   // cmd_xbar_demux:src6_data -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:cp_data
	wire   [6:0] cmd_xbar_demux_src6_channel;                                                                                // cmd_xbar_demux:src6_channel -> qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                            // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                                  // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                          // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [86:0] rsp_xbar_demux_src0_data;                                                                                   // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [6:0] rsp_xbar_demux_src0_channel;                                                                                // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                                  // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                        // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                              // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                                      // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [86:0] rsp_xbar_demux_001_src0_data;                                                                               // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [6:0] rsp_xbar_demux_001_src0_channel;                                                                            // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                              // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                        // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                              // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                                      // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [86:0] rsp_xbar_demux_002_src0_data;                                                                               // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [6:0] rsp_xbar_demux_002_src0_channel;                                                                            // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                              // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                        // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                              // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                                      // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [86:0] rsp_xbar_demux_003_src0_data;                                                                               // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [6:0] rsp_xbar_demux_003_src0_channel;                                                                            // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                              // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                        // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                              // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                                      // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [86:0] rsp_xbar_demux_004_src0_data;                                                                               // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [6:0] rsp_xbar_demux_004_src0_channel;                                                                            // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                              // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                        // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                              // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                                      // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [86:0] rsp_xbar_demux_005_src0_data;                                                                               // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [6:0] rsp_xbar_demux_005_src0_channel;                                                                            // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                              // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                        // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                              // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                                      // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [86:0] rsp_xbar_demux_006_src0_data;                                                                               // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire   [6:0] rsp_xbar_demux_006_src0_channel;                                                                            // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                              // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                                // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                              // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [86:0] limiter_cmd_src_data;                                                                                       // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [6:0] limiter_cmd_src_channel;                                                                                    // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                                      // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                               // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                                     // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                             // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [86:0] rsp_xbar_mux_src_data;                                                                                      // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [6:0] rsp_xbar_mux_src_channel;                                                                                   // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                                     // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         cmd_xbar_demux_src0_ready;                                                                                  // RGB_LED_F0_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire         id_router_src_endofpacket;                                                                                  // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                        // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                                // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [86:0] id_router_src_data;                                                                                         // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [6:0] id_router_src_channel;                                                                                      // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                        // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_demux_src1_ready;                                                                                  // RGB_LED_F1_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire         id_router_001_src_endofpacket;                                                                              // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                                    // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                            // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [86:0] id_router_001_src_data;                                                                                     // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [6:0] id_router_001_src_channel;                                                                                  // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                                    // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_src2_ready;                                                                                  // RGB_LED_F2_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	wire         id_router_002_src_endofpacket;                                                                              // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                                    // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                            // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [86:0] id_router_002_src_data;                                                                                     // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [6:0] id_router_002_src_channel;                                                                                  // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                                    // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_src3_ready;                                                                                  // RGB_LED_F3_LEDD_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src3_ready
	wire         id_router_003_src_endofpacket;                                                                              // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                                    // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                            // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [86:0] id_router_003_src_data;                                                                                     // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [6:0] id_router_003_src_channel;                                                                                  // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                                    // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_src4_ready;                                                                                  // TEST_REG_0_TestReg_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src4_ready
	wire         id_router_004_src_endofpacket;                                                                              // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                                    // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                            // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [86:0] id_router_004_src_data;                                                                                     // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [6:0] id_router_004_src_channel;                                                                                  // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                                    // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_src5_ready;                                                                                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src5_ready
	wire         id_router_005_src_endofpacket;                                                                              // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                                    // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                            // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [86:0] id_router_005_src_data;                                                                                     // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [6:0] id_router_005_src_channel;                                                                                  // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                                    // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_src6_ready;                                                                                  // qsys_basic_lophilo_module_ctrl_0_Ctrl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src6_ready
	wire         id_router_006_src_endofpacket;                                                                              // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                                    // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                            // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [86:0] id_router_006_src_data;                                                                                     // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [6:0] id_router_006_src_channel;                                                                                  // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                                    // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire   [6:0] limiter_cmd_valid_data;                                                                                     // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                                   // qsys_basic_lophilo_module_ctrl_0:ins_OC_irq -> irq_mapper:receiver0_irq
	wire   [9:0] sam9_host_events_irq;                                                                                       // irq_synchronizer:sender_irq -> SAM9_HOST:inr_EVENTS_irq
	wire   [9:0] irq_synchronizer_receiver_irq;                                                                              // irq_mapper:sender_irq -> irq_synchronizer:receiver_irq

	qsys_host_SAM9 sam9_host (
		.rso_MRST_reset       (sam9_host_mrst_reset),       //   MRST.reset
		.cso_MCLK_clk         (sam9_host_mclk_clk),         //   MCLK.clk
		.cso_H1CLK_clk        (),                           //  H1CLK.clk
		.cso_H2CLK_clk        (),                           //  H2CLK.clk
		.avm_M1_writedata     (sam9_host_m1_writedata),     //     M1.writedata
		.avm_M1_readdata      (sam9_host_m1_readdata),      //       .readdata
		.avm_M1_address       (sam9_host_m1_address),       //       .address
		.avm_M1_byteenable    (sam9_host_m1_byteenable),    //       .byteenable
		.avm_M1_write         (sam9_host_m1_write),         //       .write
		.avm_M1_read          (sam9_host_m1_read),          //       .read
		.avm_M1_begintransfer (sam9_host_m1_begintransfer), //       .begintransfer
		.avm_M1_readdatavalid (sam9_host_m1_readdatavalid), //       .readdatavalid
		.avm_M1_waitrequest   (sam9_host_m1_waitrequest),   //       .waitrequest
		.inr_EVENTS_irq       (sam9_host_events_irq),       // EVENTS.irq
		.coe_M1_RSTN          (m1_RSTN),                    // EXPORT.export
		.coe_M1_CLK           (m1_CLK),                     //       .export
		.coe_M1_ADDR          (m1_ADDR),                    //       .export
		.coe_M1_DATA          (m1_DATA),                    //       .export
		.coe_M1_CSN           (m1_CSN),                     //       .export
		.coe_M1_BEN           (m1_BEN),                     //       .export
		.coe_M1_RDN           (m1_RDN),                     //       .export
		.coe_M1_WRN           (m1_WRN),                     //       .export
		.coe_M1_WAITN         (m1_WAITN),                   //       .export
		.coe_M1_EINT          (m1_EINT)                     //       .export
	);

	qsys_basic_RGB_LED rgb_led_f0 (
		.rsi_MRST_reset       (sam9_host_mrst_reset),                                       //   MRST.reset
		.csi_MCLK_clk         (sam9_host_mclk_clk),                                         //   MCLK.clk
		.avs_LEDD_writedata   (rgb_led_f0_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (rgb_led_f0_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (rgb_led_f0_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (rgb_led_f0_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (rgb_led_f0_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (rgb_led_f0_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (rgb_led_f0s_leds_data),                                      //   LEDS.data
		.asi_LEDS_valid       (rgb_led_f0s_leds_valid),                                     //       .valid
		.asi_LEDS_ready       (rgb_led_f0s_leds_ready),                                     //       .ready
		.coe_LED_R            (led_f0_R),                                                   // EXPORT.export
		.coe_LED_G            (led_f0_G),                                                   //       .export
		.coe_LED_B            (led_f0_B)                                                    //       .export
	);

	qsys_basic_RGB_LED rgb_led_f1 (
		.rsi_MRST_reset       (sam9_host_mrst_reset),                                       //   MRST.reset
		.csi_MCLK_clk         (sam9_host_mclk_clk),                                         //   MCLK.clk
		.avs_LEDD_writedata   (rgb_led_f1_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (rgb_led_f1_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (rgb_led_f1_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (rgb_led_f1_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (rgb_led_f1_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (rgb_led_f1_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (rgb_led_f1s_leds_data),                                      //   LEDS.data
		.asi_LEDS_valid       (rgb_led_f1s_leds_valid),                                     //       .valid
		.asi_LEDS_ready       (rgb_led_f1s_leds_ready),                                     //       .ready
		.coe_LED_R            (led_f1_R),                                                   // EXPORT.export
		.coe_LED_G            (led_f1_G),                                                   //       .export
		.coe_LED_B            (led_f1_B)                                                    //       .export
	);

	qsys_basic_RGB_LED rgb_led_f2 (
		.rsi_MRST_reset       (sam9_host_mrst_reset),                                       //   MRST.reset
		.csi_MCLK_clk         (sam9_host_mclk_clk),                                         //   MCLK.clk
		.avs_LEDD_writedata   (rgb_led_f2_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (rgb_led_f2_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (rgb_led_f2_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (rgb_led_f2_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (rgb_led_f2_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (rgb_led_f2_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (rgb_led_f2s_leds_data),                                      //   LEDS.data
		.asi_LEDS_valid       (rgb_led_f2s_leds_valid),                                     //       .valid
		.asi_LEDS_ready       (rgb_led_f2s_leds_ready),                                     //       .ready
		.coe_LED_R            (led_f2_R),                                                   // EXPORT.export
		.coe_LED_G            (led_f2_G),                                                   //       .export
		.coe_LED_B            (led_f2_B)                                                    //       .export
	);

	qsys_basic_RGB_LED rgb_led_f3 (
		.rsi_MRST_reset       (sam9_host_mrst_reset),                                       //   MRST.reset
		.csi_MCLK_clk         (sam9_host_mclk_clk),                                         //   MCLK.clk
		.avs_LEDD_writedata   (rgb_led_f3_ledd_translator_avalon_anti_slave_0_writedata),   //   LEDD.writedata
		.avs_LEDD_readdata    (rgb_led_f3_ledd_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_LEDD_byteenable  (rgb_led_f3_ledd_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_LEDD_write       (rgb_led_f3_ledd_translator_avalon_anti_slave_0_write),       //       .write
		.avs_LEDD_read        (rgb_led_f3_ledd_translator_avalon_anti_slave_0_read),        //       .read
		.avs_LEDD_waitrequest (rgb_led_f3_ledd_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.asi_LEDS_data        (rgb_led_f3s_leds_data),                                      //   LEDS.data
		.asi_LEDS_valid       (rgb_led_f3s_leds_valid),                                     //       .valid
		.asi_LEDS_ready       (rgb_led_f3s_leds_ready),                                     //       .ready
		.coe_LED_R            (led_f3_R),                                                   // EXPORT.export
		.coe_LED_G            (led_f3_G),                                                   //       .export
		.coe_LED_B            (led_f3_B)                                                    //       .export
	);

	qsys_test_RGB_LED_ASO rgb_led_f0s (
		.rsi_MRST_reset (sam9_host_mrst_reset),   // MRST.reset
		.csi_MCLK_clk   (sam9_host_mclk_clk),     // MCLK.clk
		.aso_LEDS_data  (rgb_led_f0s_leds_data),  // LEDS.data
		.aso_LEDS_valid (rgb_led_f0s_leds_valid), //     .valid
		.aso_LEDS_ready (rgb_led_f0s_leds_ready)  //     .ready
	);

	qsys_test_RGB_LED_ASO rgb_led_f1s (
		.rsi_MRST_reset (sam9_host_mrst_reset),   // MRST.reset
		.csi_MCLK_clk   (sam9_host_mclk_clk),     // MCLK.clk
		.aso_LEDS_data  (rgb_led_f1s_leds_data),  // LEDS.data
		.aso_LEDS_valid (rgb_led_f1s_leds_valid), //     .valid
		.aso_LEDS_ready (rgb_led_f1s_leds_ready)  //     .ready
	);

	qsys_test_RGB_LED_ASO rgb_led_f2s (
		.rsi_MRST_reset (sam9_host_mrst_reset),   // MRST.reset
		.csi_MCLK_clk   (sam9_host_mclk_clk),     // MCLK.clk
		.aso_LEDS_data  (rgb_led_f2s_leds_data),  // LEDS.data
		.aso_LEDS_valid (rgb_led_f2s_leds_valid), //     .valid
		.aso_LEDS_ready (rgb_led_f2s_leds_ready)  //     .ready
	);

	qsys_test_RGB_LED_ASO rgb_led_f3s (
		.rsi_MRST_reset (sam9_host_mrst_reset),   // MRST.reset
		.csi_MCLK_clk   (sam9_host_mclk_clk),     // MCLK.clk
		.aso_LEDS_data  (rgb_led_f3s_leds_data),  // LEDS.data
		.aso_LEDS_valid (rgb_led_f3s_leds_valid), //     .valid
		.aso_LEDS_ready (rgb_led_f3s_leds_ready)  //     .ready
	);

	qsys_test_RegRW test_reg_0 (
		.rsi_MRST_reset          (sam9_host_mrst_reset),                                          //    MRST.reset
		.csi_MCLK_clk            (sam9_host_mclk_clk),                                            //    MCLK.clk
		.avs_TestReg_readdata    (test_reg_0_testreg_translator_avalon_anti_slave_0_readdata),    // TestReg.readdata
		.avs_TestReg_read        (test_reg_0_testreg_translator_avalon_anti_slave_0_read),        //        .read
		.avs_TestReg_writedata   (test_reg_0_testreg_translator_avalon_anti_slave_0_writedata),   //        .writedata
		.avs_TestReg_write       (test_reg_0_testreg_translator_avalon_anti_slave_0_write),       //        .write
		.avs_TestReg_waitrequest (test_reg_0_testreg_translator_avalon_anti_slave_0_waitrequest)  //        .waitrequest
	);

	frontier_onchip_memory2_0 onchip_memory2_0 (
		.clk        (sam9_host_mclk_clk),                                            //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (sam9_host_mrst_reset)                                           // reset1.reset
	);

	qsys_basic_lophilo_module_ctrl qsys_basic_lophilo_module_ctrl_0 (
		.rsi_MRST_reset       (sam9_host_mrst_reset),                                                             //   MRST.reset
		.csi_MCLK_clk         (sam9_host_mclk_clk),                                                               //   MCLK.clk
		.avs_Ctrl_writedata   (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_writedata),   //   Ctrl.writedata
		.avs_Ctrl_readdata    (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_readdata),    //       .readdata
		.avs_Ctrl_byteenable  (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_byteenable),  //       .byteenable
		.avs_Ctrl_write       (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_write),       //       .write
		.avs_Ctrl_read        (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_read),        //       .read
		.avs_Ctrl_waitrequest (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_waitrequest), //       .waitrequest
		.ins_OC_irq           (irq_mapper_receiver0_irq),                                                         //     OC.irq
		.coe_A_OCN            (admin_A_OCN),                                                                      // EXPORT.export
		.coe_A_PWREN          (admin_A_PWREN),                                                                    //       .export
		.coe_A_HOE            (admin_A_HOE),                                                                      //       .export
		.coe_A_LOE            (admin_A_LOE),                                                                      //       .export
		.coe_B_OCN            (admin_B_OCN),                                                                      //       .export
		.coe_B_PWREN          (admin_B_PWREN),                                                                    //       .export
		.coe_B_HOE            (admin_B_HOE),                                                                      //       .export
		.coe_B_LOE            (admin_B_LOE)                                                                       //       .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (1),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sam9_host_m1_translator (
		.clk                   (sam9_host_mclk_clk),                                              //                       clk.clk
		.reset                 (sam9_host_mrst_reset),                                            //                     reset.reset
		.uav_address           (sam9_host_m1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sam9_host_m1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sam9_host_m1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sam9_host_m1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sam9_host_m1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sam9_host_m1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sam9_host_m1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sam9_host_m1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sam9_host_m1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sam9_host_m1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sam9_host_m1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sam9_host_m1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sam9_host_m1_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (sam9_host_m1_byteenable),                                         //                          .byteenable
		.av_begintransfer      (sam9_host_m1_begintransfer),                                      //                          .begintransfer
		.av_read               (sam9_host_m1_read),                                               //                          .read
		.av_readdata           (sam9_host_m1_readdata),                                           //                          .readdata
		.av_readdatavalid      (sam9_host_m1_readdatavalid),                                      //                          .readdatavalid
		.av_write              (sam9_host_m1_write),                                              //                          .write
		.av_writedata          (sam9_host_m1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                            //               (terminated)
		.av_chipselect         (1'b0),                                                            //               (terminated)
		.av_lock               (1'b0),                                                            //               (terminated)
		.av_debugaccess        (1'b0),                                                            //               (terminated)
		.uav_clken             (),                                                                //               (terminated)
		.av_clken              (1'b1)                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rgb_led_f0_ledd_translator (
		.clk                   (sam9_host_mclk_clk),                                                         //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                       //                    reset.reset
		.uav_address           (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (rgb_led_f0_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (rgb_led_f0_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (rgb_led_f0_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (rgb_led_f0_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (rgb_led_f0_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (rgb_led_f0_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                           //              (terminated)
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_burstcount         (),                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_lock               (),                                                                           //              (terminated)
		.av_chipselect         (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_debugaccess        (),                                                                           //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rgb_led_f1_ledd_translator (
		.clk                   (sam9_host_mclk_clk),                                                         //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                       //                    reset.reset
		.uav_address           (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (rgb_led_f1_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (rgb_led_f1_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (rgb_led_f1_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (rgb_led_f1_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (rgb_led_f1_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (rgb_led_f1_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                           //              (terminated)
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_burstcount         (),                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_lock               (),                                                                           //              (terminated)
		.av_chipselect         (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_debugaccess        (),                                                                           //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rgb_led_f2_ledd_translator (
		.clk                   (sam9_host_mclk_clk),                                                         //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                       //                    reset.reset
		.uav_address           (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (rgb_led_f2_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (rgb_led_f2_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (rgb_led_f2_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (rgb_led_f2_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (rgb_led_f2_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (rgb_led_f2_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                           //              (terminated)
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_burstcount         (),                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_lock               (),                                                                           //              (terminated)
		.av_chipselect         (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_debugaccess        (),                                                                           //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rgb_led_f3_ledd_translator (
		.clk                   (sam9_host_mclk_clk),                                                         //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                       //                    reset.reset
		.uav_address           (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (rgb_led_f3_ledd_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (rgb_led_f3_ledd_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (rgb_led_f3_ledd_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (rgb_led_f3_ledd_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (rgb_led_f3_ledd_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (rgb_led_f3_ledd_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                           //              (terminated)
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_burstcount         (),                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_lock               (),                                                                           //              (terminated)
		.av_chipselect         (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_debugaccess        (),                                                                           //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) test_reg_0_testreg_translator (
		.clk                   (sam9_host_mclk_clk),                                                            //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                          //                    reset.reset
		.uav_address           (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (test_reg_0_testreg_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (test_reg_0_testreg_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (test_reg_0_testreg_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (test_reg_0_testreg_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (test_reg_0_testreg_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                   (sam9_host_mclk_clk),                                                             //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                           //                    reset.reset
		.uav_address           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) qsys_basic_lophilo_module_ctrl_0_ctrl_translator (
		.clk                   (sam9_host_mclk_clk),                                                                               //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                                             //                    reset.reset
		.uav_address           (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                                                 //              (terminated)
		.av_begintransfer      (),                                                                                                 //              (terminated)
		.av_beginbursttransfer (),                                                                                                 //              (terminated)
		.av_burstcount         (),                                                                                                 //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable    (),                                                                                                 //              (terminated)
		.av_lock               (),                                                                                                 //              (terminated)
		.av_chipselect         (),                                                                                                 //              (terminated)
		.av_clken              (),                                                                                                 //              (terminated)
		.uav_clken             (1'b0),                                                                                             //              (terminated)
		.av_debugaccess        (),                                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                                  //              (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                                   //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                                 //       clk_reset.reset
		.m0_address              (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src2_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_src2_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_src2_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_src2_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src2_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src2_channel),                                                          //                .channel
		.rf_sink_ready           (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                                   //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                                 // clk_reset.reset
		.in_data           (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                                   //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                                 //       clk_reset.reset
		.m0_address              (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src3_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_src3_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_src3_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_src3_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src3_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src3_channel),                                                          //                .channel
		.rf_sink_ready           (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                                   //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                                 // clk_reset.reset
		.in_data           (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                                   //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                                 //       clk_reset.reset
		.m0_address              (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                          //                .channel
		.rf_sink_ready           (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                                   //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                                 // clk_reset.reset
		.in_data           (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) test_reg_0_testreg_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                                      //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                                    //       clk_reset.reset
		.m0_address              (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src4_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_src4_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_src4_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_src4_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src4_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src4_channel),                                                             //                .channel
		.rf_sink_ready           (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                                      //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                                    // clk_reset.reset
		.in_data           (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                                   //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                                 //       clk_reset.reset
		.m0_address              (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                          //                .channel
		.rf_sink_ready           (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                                   //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                                 // clk_reset.reset
		.in_data           (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (7),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7)
	) sam9_host_m1_translator_avalon_universal_master_0_agent (
		.clk              (sam9_host_mclk_clk),                                                       //       clk.clk
		.reset            (sam9_host_mrst_reset),                                                     // clk_reset.reset
		.av_address       (sam9_host_m1_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sam9_host_m1_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sam9_host_m1_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sam9_host_m1_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sam9_host_m1_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sam9_host_m1_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sam9_host_m1_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sam9_host_m1_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sam9_host_m1_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sam9_host_m1_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sam9_host_m1_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                    //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                     //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                  //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                     //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                                       //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                                     //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src5_ready),                                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_src5_valid),                                                                //                .valid
		.cp_data                 (cmd_xbar_demux_src5_data),                                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_src5_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src5_endofpacket),                                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src5_channel),                                                              //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                                       //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                                     // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (7),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                                                         //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                                                       //       clk_reset.reset
		.m0_address              (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src6_ready),                                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_src6_valid),                                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_src6_data),                                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_src6_startofpacket),                                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src6_endofpacket),                                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src6_channel),                                                                                //                .channel
		.rf_sink_ready           (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                                                         //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                                                       // clk_reset.reset
		.in_data           (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	frontier_addr_router addr_router (
		.sink_ready         (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                       //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_src_valid),                                                    //          .valid
		.src_data           (addr_router_src_data),                                                     //          .data
		.src_channel        (addr_router_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                               //          .endofpacket
	);

	frontier_id_router id_router (
		.sink_ready         (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rgb_led_f0_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                         //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                        //       src.ready
		.src_valid          (id_router_src_valid),                                                        //          .valid
		.src_data           (id_router_src_data),                                                         //          .data
		.src_channel        (id_router_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                   //          .endofpacket
	);

	frontier_id_router id_router_001 (
		.sink_ready         (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rgb_led_f1_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                         //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                    //       src.ready
		.src_valid          (id_router_001_src_valid),                                                    //          .valid
		.src_data           (id_router_001_src_data),                                                     //          .data
		.src_channel        (id_router_001_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                               //          .endofpacket
	);

	frontier_id_router id_router_002 (
		.sink_ready         (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rgb_led_f2_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                         //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                    //       src.ready
		.src_valid          (id_router_002_src_valid),                                                    //          .valid
		.src_data           (id_router_002_src_data),                                                     //          .data
		.src_channel        (id_router_002_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                               //          .endofpacket
	);

	frontier_id_router id_router_003 (
		.sink_ready         (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rgb_led_f3_ledd_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                         //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                    //       src.ready
		.src_valid          (id_router_003_src_valid),                                                    //          .valid
		.src_data           (id_router_003_src_data),                                                     //          .data
		.src_channel        (id_router_003_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                               //          .endofpacket
	);

	frontier_id_router id_router_004 (
		.sink_ready         (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (test_reg_0_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                            //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                       //       src.ready
		.src_valid          (id_router_004_src_valid),                                                       //          .valid
		.src_data           (id_router_004_src_data),                                                        //          .data
		.src_channel        (id_router_004_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                  //          .endofpacket
	);

	frontier_id_router id_router_005 (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                             //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                        //       src.ready
		.src_valid          (id_router_005_src_valid),                                                        //          .valid
		.src_data           (id_router_005_src_data),                                                         //          .data
		.src_channel        (id_router_005_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                   //          .endofpacket
	);

	frontier_id_router id_router_006 (
		.sink_ready         (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (qsys_basic_lophilo_module_ctrl_0_ctrl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                                               //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                                             // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                          //          .valid
		.src_data           (id_router_006_src_data),                                                                           //          .data
		.src_channel        (id_router_006_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                                     //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (7),
		.VALID_WIDTH               (7),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (sam9_host_mclk_clk),             //       clk.clk
		.reset                  (sam9_host_mrst_reset),           // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	frontier_cmd_xbar_demux cmd_xbar_demux (
		.clk                (sam9_host_mclk_clk),                //        clk.clk
		.reset              (sam9_host_mrst_reset),              //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_src6_endofpacket)    //           .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux (
		.clk                (sam9_host_mclk_clk),                //       clk.clk
		.reset              (sam9_host_mrst_reset),              // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (sam9_host_mclk_clk),                    //       clk.clk
		.reset              (sam9_host_mrst_reset),                  // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (sam9_host_mclk_clk),                    //       clk.clk
		.reset              (sam9_host_mrst_reset),                  // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (sam9_host_mclk_clk),                    //       clk.clk
		.reset              (sam9_host_mrst_reset),                  // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (sam9_host_mclk_clk),                    //       clk.clk
		.reset              (sam9_host_mrst_reset),                  // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (sam9_host_mclk_clk),                    //       clk.clk
		.reset              (sam9_host_mrst_reset),                  // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (sam9_host_mclk_clk),                    //       clk.clk
		.reset              (sam9_host_mrst_reset),                  // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (sam9_host_mclk_clk),                    //       clk.clk
		.reset               (sam9_host_mrst_reset),                  // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	frontier_irq_mapper irq_mapper (
		.clk           (sam9_host_mclk_clk),            //       clk.clk
		.reset         (sam9_host_mrst_reset),          // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),      // receiver0.irq
		.sender_irq    (irq_synchronizer_receiver_irq)  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (10)
	) irq_synchronizer (
		.receiver_clk   (sam9_host_mclk_clk),            //       receiver_clk.clk
		.sender_clk     (sam9_host_mclk_clk),            //         sender_clk.clk
		.receiver_reset (sam9_host_mrst_reset),          // receiver_clk_reset.reset
		.sender_reset   (sam9_host_mrst_reset),          //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq), //           receiver.irq
		.sender_irq     (sam9_host_events_irq)           //             sender.irq
	);

endmodule
