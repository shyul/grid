// frontier.v

// Generated using ACDS version 11.1sp2 259 at 2012.07.17.11:15:56

`timescale 1 ps / 1 ps
module frontier (
		output wire        led_F0R,  // led.F0R
		output wire        led_F0G,  //    .F0G
		output wire        led_F0B,  //    .F0B
		output wire        led_F1R,  //    .F1R
		output wire        led_F1G,  //    .F1G
		output wire        led_F1B,  //    .F1B
		output wire        led_F2R,  //    .F2R
		output wire        led_F2G,  //    .F2G
		output wire        led_F2B,  //    .F2B
		output wire        led_F3R,  //    .F3R
		output wire        led_F3G,  //    .F3G
		output wire        led_F3B,  //    .F3B
		input  wire        m1_RSTN,  //  m1.RSTN
		input  wire        m1_CLK,   //    .CLK
		input  wire [21:0] m1_ADDR,  //    .ADDR
		inout  wire [31:0] m1_DATA,  //    .DATA
		input  wire [3:0]  m1_CSN,   //    .CSN
		input  wire [3:0]  m1_BEN,   //    .BEN
		input  wire        m1_RDN,   //    .RDN
		input  wire        m1_WRN,   //    .WRN
		output wire        m1_WAITN, //    .WAITN
		output wire [9:0]  m1_EINT   //    .EINT
	);

	wire         sam9_host_mrst_reset;                                                                   // SAM9_HOST:rso_MRST_reset -> [SAM9_HOST_M1_translator:reset, SAM9_HOST_M1_translator_avalon_universal_master_0_agent:reset, TEST_LED:rsi_MRST_reset, TEST_LED_TestReg_translator:reset, TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:reset, TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, TEST_MEM:reset, TEST_MEM_s1_translator:reset, TEST_MEM_s1_translator_avalon_universal_slave_0_agent:reset, TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, TEST_REG0:rsi_MRST_reset, TEST_REG0_TestReg_translator:reset, TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:reset, TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, TEST_REG1:rsi_MRST_reset, TEST_REG1_TestReg_translator:reset, TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:reset, TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, TEST_REG2:rsi_MRST_reset, TEST_REG2_TestReg_translator:reset, TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:reset, TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, cmd_xbar_demux:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, irq_mapper:reset, irq_synchronizer:receiver_reset, irq_synchronizer:sender_reset, limiter:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_mux:reset]
	wire         sam9_host_mclk_clk;                                                                     // SAM9_HOST:cso_MCLK_clk -> [SAM9_HOST_M1_translator:clk, SAM9_HOST_M1_translator_avalon_universal_master_0_agent:clk, TEST_LED:csi_MCLK_clk, TEST_LED_TestReg_translator:clk, TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:clk, TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, TEST_MEM:clk, TEST_MEM_s1_translator:clk, TEST_MEM_s1_translator_avalon_universal_slave_0_agent:clk, TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, TEST_REG0:csi_MCLK_clk, TEST_REG0_TestReg_translator:clk, TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:clk, TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, TEST_REG1:csi_MCLK_clk, TEST_REG1_TestReg_translator:clk, TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:clk, TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, TEST_REG2:csi_MCLK_clk, TEST_REG2_TestReg_translator:clk, TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:clk, TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, cmd_xbar_demux:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, irq_mapper:clk, irq_synchronizer:receiver_clk, irq_synchronizer:sender_clk, limiter:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_mux:clk]
	wire         sam9_host_m1_waitrequest;                                                               // SAM9_HOST_M1_translator:av_waitrequest -> SAM9_HOST:avm_M1_waitrequest
	wire  [31:0] sam9_host_m1_address;                                                                   // SAM9_HOST:avm_M1_address -> SAM9_HOST_M1_translator:av_address
	wire  [31:0] sam9_host_m1_writedata;                                                                 // SAM9_HOST:avm_M1_writedata -> SAM9_HOST_M1_translator:av_writedata
	wire         sam9_host_m1_write;                                                                     // SAM9_HOST:avm_M1_write -> SAM9_HOST_M1_translator:av_write
	wire         sam9_host_m1_read;                                                                      // SAM9_HOST:avm_M1_read -> SAM9_HOST_M1_translator:av_read
	wire  [31:0] sam9_host_m1_readdata;                                                                  // SAM9_HOST_M1_translator:av_readdata -> SAM9_HOST:avm_M1_readdata
	wire         sam9_host_m1_begintransfer;                                                             // SAM9_HOST:avm_M1_begintransfer -> SAM9_HOST_M1_translator:av_begintransfer
	wire         sam9_host_m1_readdatavalid;                                                             // SAM9_HOST_M1_translator:av_readdatavalid -> SAM9_HOST:avm_M1_readdatavalid
	wire   [3:0] sam9_host_m1_byteenable;                                                                // SAM9_HOST:avm_M1_byteenable -> SAM9_HOST_M1_translator:av_byteenable
	wire         test_led_testreg_translator_avalon_anti_slave_0_waitrequest;                            // TEST_LED:avs_TestReg_waitrequest -> TEST_LED_TestReg_translator:av_waitrequest
	wire  [31:0] test_led_testreg_translator_avalon_anti_slave_0_writedata;                              // TEST_LED_TestReg_translator:av_writedata -> TEST_LED:avs_TestReg_writedata
	wire         test_led_testreg_translator_avalon_anti_slave_0_write;                                  // TEST_LED_TestReg_translator:av_write -> TEST_LED:avs_TestReg_write
	wire         test_led_testreg_translator_avalon_anti_slave_0_read;                                   // TEST_LED_TestReg_translator:av_read -> TEST_LED:avs_TestReg_read
	wire  [31:0] test_led_testreg_translator_avalon_anti_slave_0_readdata;                               // TEST_LED:avs_TestReg_readdata -> TEST_LED_TestReg_translator:av_readdata
	wire         test_reg0_testreg_translator_avalon_anti_slave_0_waitrequest;                           // TEST_REG0:avs_TestReg_waitrequest -> TEST_REG0_TestReg_translator:av_waitrequest
	wire  [31:0] test_reg0_testreg_translator_avalon_anti_slave_0_writedata;                             // TEST_REG0_TestReg_translator:av_writedata -> TEST_REG0:avs_TestReg_writedata
	wire         test_reg0_testreg_translator_avalon_anti_slave_0_write;                                 // TEST_REG0_TestReg_translator:av_write -> TEST_REG0:avs_TestReg_write
	wire         test_reg0_testreg_translator_avalon_anti_slave_0_read;                                  // TEST_REG0_TestReg_translator:av_read -> TEST_REG0:avs_TestReg_read
	wire  [31:0] test_reg0_testreg_translator_avalon_anti_slave_0_readdata;                              // TEST_REG0:avs_TestReg_readdata -> TEST_REG0_TestReg_translator:av_readdata
	wire         test_reg1_testreg_translator_avalon_anti_slave_0_waitrequest;                           // TEST_REG1:avs_TestReg_waitrequest -> TEST_REG1_TestReg_translator:av_waitrequest
	wire  [31:0] test_reg1_testreg_translator_avalon_anti_slave_0_writedata;                             // TEST_REG1_TestReg_translator:av_writedata -> TEST_REG1:avs_TestReg_writedata
	wire         test_reg1_testreg_translator_avalon_anti_slave_0_write;                                 // TEST_REG1_TestReg_translator:av_write -> TEST_REG1:avs_TestReg_write
	wire         test_reg1_testreg_translator_avalon_anti_slave_0_read;                                  // TEST_REG1_TestReg_translator:av_read -> TEST_REG1:avs_TestReg_read
	wire  [31:0] test_reg1_testreg_translator_avalon_anti_slave_0_readdata;                              // TEST_REG1:avs_TestReg_readdata -> TEST_REG1_TestReg_translator:av_readdata
	wire         test_reg2_testreg_translator_avalon_anti_slave_0_waitrequest;                           // TEST_REG2:avs_TestReg_waitrequest -> TEST_REG2_TestReg_translator:av_waitrequest
	wire  [31:0] test_reg2_testreg_translator_avalon_anti_slave_0_writedata;                             // TEST_REG2_TestReg_translator:av_writedata -> TEST_REG2:avs_TestReg_writedata
	wire         test_reg2_testreg_translator_avalon_anti_slave_0_write;                                 // TEST_REG2_TestReg_translator:av_write -> TEST_REG2:avs_TestReg_write
	wire         test_reg2_testreg_translator_avalon_anti_slave_0_read;                                  // TEST_REG2_TestReg_translator:av_read -> TEST_REG2:avs_TestReg_read
	wire  [31:0] test_reg2_testreg_translator_avalon_anti_slave_0_readdata;                              // TEST_REG2:avs_TestReg_readdata -> TEST_REG2_TestReg_translator:av_readdata
	wire  [31:0] test_mem_s1_translator_avalon_anti_slave_0_writedata;                                   // TEST_MEM_s1_translator:av_writedata -> TEST_MEM:writedata
	wire   [9:0] test_mem_s1_translator_avalon_anti_slave_0_address;                                     // TEST_MEM_s1_translator:av_address -> TEST_MEM:address
	wire         test_mem_s1_translator_avalon_anti_slave_0_chipselect;                                  // TEST_MEM_s1_translator:av_chipselect -> TEST_MEM:chipselect
	wire         test_mem_s1_translator_avalon_anti_slave_0_clken;                                       // TEST_MEM_s1_translator:av_clken -> TEST_MEM:clken
	wire         test_mem_s1_translator_avalon_anti_slave_0_write;                                       // TEST_MEM_s1_translator:av_write -> TEST_MEM:write
	wire  [31:0] test_mem_s1_translator_avalon_anti_slave_0_readdata;                                    // TEST_MEM:readdata -> TEST_MEM_s1_translator:av_readdata
	wire   [3:0] test_mem_s1_translator_avalon_anti_slave_0_byteenable;                                  // TEST_MEM_s1_translator:av_byteenable -> TEST_MEM:byteenable
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // TEST_REG2_TestReg_translator:uav_waitrequest -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount;              // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:m0_burstcount -> TEST_REG2_TestReg_translator:uav_burstcount
	wire  [31:0] test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_writedata;               // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:m0_writedata -> TEST_REG2_TestReg_translator:uav_writedata
	wire  [31:0] test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_address;                 // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:m0_address -> TEST_REG2_TestReg_translator:uav_address
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_write;                   // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:m0_write -> TEST_REG2_TestReg_translator:uav_write
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_lock;                    // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:m0_lock -> TEST_REG2_TestReg_translator:uav_lock
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_read;                    // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:m0_read -> TEST_REG2_TestReg_translator:uav_read
	wire  [31:0] test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_readdata;                // TEST_REG2_TestReg_translator:uav_readdata -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // TEST_REG2_TestReg_translator:uav_readdatavalid -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:m0_debugaccess -> TEST_REG2_TestReg_translator:uav_debugaccess
	wire   [3:0] test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable;              // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:m0_byteenable -> TEST_REG2_TestReg_translator:uav_byteenable
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid;            // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rf_source_valid -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_data;             // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rf_source_data -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready;            // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_ready -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] test_reg2_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // TEST_MEM_s1_translator:uav_waitrequest -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] test_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> TEST_MEM_s1_translator:uav_burstcount
	wire  [31:0] test_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                     // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> TEST_MEM_s1_translator:uav_writedata
	wire  [31:0] test_mem_s1_translator_avalon_universal_slave_0_agent_m0_address;                       // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:m0_address -> TEST_MEM_s1_translator:uav_address
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_m0_write;                         // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:m0_write -> TEST_MEM_s1_translator:uav_write
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock;                          // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> TEST_MEM_s1_translator:uav_lock
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_m0_read;                          // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:m0_read -> TEST_MEM_s1_translator:uav_read
	wire  [31:0] test_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                      // TEST_MEM_s1_translator:uav_readdata -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // TEST_MEM_s1_translator:uav_readdatavalid -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> TEST_MEM_s1_translator:uav_debugaccess
	wire   [3:0] test_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> TEST_MEM_s1_translator:uav_byteenable
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                   // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] test_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // TEST_REG0_TestReg_translator:uav_waitrequest -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount;              // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:m0_burstcount -> TEST_REG0_TestReg_translator:uav_burstcount
	wire  [31:0] test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_writedata;               // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:m0_writedata -> TEST_REG0_TestReg_translator:uav_writedata
	wire  [31:0] test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_address;                 // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:m0_address -> TEST_REG0_TestReg_translator:uav_address
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_write;                   // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:m0_write -> TEST_REG0_TestReg_translator:uav_write
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_lock;                    // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:m0_lock -> TEST_REG0_TestReg_translator:uav_lock
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_read;                    // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:m0_read -> TEST_REG0_TestReg_translator:uav_read
	wire  [31:0] test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_readdata;                // TEST_REG0_TestReg_translator:uav_readdata -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // TEST_REG0_TestReg_translator:uav_readdatavalid -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:m0_debugaccess -> TEST_REG0_TestReg_translator:uav_debugaccess
	wire   [3:0] test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable;              // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:m0_byteenable -> TEST_REG0_TestReg_translator:uav_byteenable
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid;            // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rf_source_valid -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_data;             // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rf_source_data -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready;            // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_ready -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] test_reg0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // TEST_REG1_TestReg_translator:uav_waitrequest -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount;              // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:m0_burstcount -> TEST_REG1_TestReg_translator:uav_burstcount
	wire  [31:0] test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_writedata;               // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:m0_writedata -> TEST_REG1_TestReg_translator:uav_writedata
	wire  [31:0] test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_address;                 // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:m0_address -> TEST_REG1_TestReg_translator:uav_address
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_write;                   // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:m0_write -> TEST_REG1_TestReg_translator:uav_write
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_lock;                    // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:m0_lock -> TEST_REG1_TestReg_translator:uav_lock
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_read;                    // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:m0_read -> TEST_REG1_TestReg_translator:uav_read
	wire  [31:0] test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_readdata;                // TEST_REG1_TestReg_translator:uav_readdata -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // TEST_REG1_TestReg_translator:uav_readdatavalid -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:m0_debugaccess -> TEST_REG1_TestReg_translator:uav_debugaccess
	wire   [3:0] test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable;              // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:m0_byteenable -> TEST_REG1_TestReg_translator:uav_byteenable
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid;            // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rf_source_valid -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_data;             // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rf_source_data -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready;            // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_ready -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] test_reg1_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // TEST_LED_TestReg_translator:uav_waitrequest -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] test_led_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount;               // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:m0_burstcount -> TEST_LED_TestReg_translator:uav_burstcount
	wire  [31:0] test_led_testreg_translator_avalon_universal_slave_0_agent_m0_writedata;                // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:m0_writedata -> TEST_LED_TestReg_translator:uav_writedata
	wire  [31:0] test_led_testreg_translator_avalon_universal_slave_0_agent_m0_address;                  // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:m0_address -> TEST_LED_TestReg_translator:uav_address
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_m0_write;                    // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:m0_write -> TEST_LED_TestReg_translator:uav_write
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_m0_lock;                     // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:m0_lock -> TEST_LED_TestReg_translator:uav_lock
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_m0_read;                     // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:m0_read -> TEST_LED_TestReg_translator:uav_read
	wire  [31:0] test_led_testreg_translator_avalon_universal_slave_0_agent_m0_readdata;                 // TEST_LED_TestReg_translator:uav_readdata -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // TEST_LED_TestReg_translator:uav_readdatavalid -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:m0_debugaccess -> TEST_LED_TestReg_translator:uav_debugaccess
	wire   [3:0] test_led_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable;               // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:m0_byteenable -> TEST_LED_TestReg_translator:uav_byteenable
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid;             // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rf_source_valid -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [87:0] test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_data;              // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rf_source_data -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready;             // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [87:0] test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rf_sink_ready -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] test_led_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sam9_host_m1_translator_avalon_universal_master_0_waitrequest;                          // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_waitrequest -> SAM9_HOST_M1_translator:uav_waitrequest
	wire   [2:0] sam9_host_m1_translator_avalon_universal_master_0_burstcount;                           // SAM9_HOST_M1_translator:uav_burstcount -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] sam9_host_m1_translator_avalon_universal_master_0_writedata;                            // SAM9_HOST_M1_translator:uav_writedata -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_writedata
	wire  [31:0] sam9_host_m1_translator_avalon_universal_master_0_address;                              // SAM9_HOST_M1_translator:uav_address -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_address
	wire         sam9_host_m1_translator_avalon_universal_master_0_lock;                                 // SAM9_HOST_M1_translator:uav_lock -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_lock
	wire         sam9_host_m1_translator_avalon_universal_master_0_write;                                // SAM9_HOST_M1_translator:uav_write -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_write
	wire         sam9_host_m1_translator_avalon_universal_master_0_read;                                 // SAM9_HOST_M1_translator:uav_read -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] sam9_host_m1_translator_avalon_universal_master_0_readdata;                             // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_readdata -> SAM9_HOST_M1_translator:uav_readdata
	wire         sam9_host_m1_translator_avalon_universal_master_0_debugaccess;                          // SAM9_HOST_M1_translator:uav_debugaccess -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] sam9_host_m1_translator_avalon_universal_master_0_byteenable;                           // SAM9_HOST_M1_translator:uav_byteenable -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_byteenable
	wire         sam9_host_m1_translator_avalon_universal_master_0_readdatavalid;                        // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:av_readdatavalid -> SAM9_HOST_M1_translator:uav_readdatavalid
	wire         sam9_host_m1_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         sam9_host_m1_translator_avalon_universal_master_0_agent_cp_valid;                       // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         sam9_host_m1_translator_avalon_universal_master_0_agent_cp_startofpacket;               // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [86:0] sam9_host_m1_translator_avalon_universal_master_0_agent_cp_data;                        // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         sam9_host_m1_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router:sink_ready -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:cp_ready
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rp_valid;                    // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [86:0] test_led_testreg_translator_avalon_universal_slave_0_agent_rp_data;                     // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         test_led_testreg_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router:sink_ready -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:rp_ready
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_valid;                   // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [86:0] test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_data;                    // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_001:sink_ready -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:rp_ready
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_valid;                   // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [86:0] test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_data;                    // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_002:sink_ready -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:rp_ready
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_valid;                   // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [86:0] test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_data;                    // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_003:sink_ready -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:rp_ready
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid;                         // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [86:0] test_mem_s1_translator_avalon_universal_slave_0_agent_rp_data;                          // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         test_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_004:sink_ready -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                            // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                  // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                          // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [86:0] addr_router_src_data;                                                                   // addr_router:src_data -> limiter:cmd_sink_data
	wire   [4:0] addr_router_src_channel;                                                                // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                  // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                            // limiter:rsp_src_endofpacket -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                  // limiter:rsp_src_valid -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                          // limiter:rsp_src_startofpacket -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [86:0] limiter_rsp_src_data;                                                                   // limiter:rsp_src_data -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_data
	wire   [4:0] limiter_rsp_src_channel;                                                                // limiter:rsp_src_channel -> SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                  // SAM9_HOST_M1_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         cmd_xbar_demux_src0_endofpacket;                                                        // cmd_xbar_demux:src0_endofpacket -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                              // cmd_xbar_demux:src0_valid -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                      // cmd_xbar_demux:src0_startofpacket -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src0_data;                                                               // cmd_xbar_demux:src0_data -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:cp_data
	wire   [4:0] cmd_xbar_demux_src0_channel;                                                            // cmd_xbar_demux:src0_channel -> TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src1_endofpacket;                                                        // cmd_xbar_demux:src1_endofpacket -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                              // cmd_xbar_demux:src1_valid -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                      // cmd_xbar_demux:src1_startofpacket -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src1_data;                                                               // cmd_xbar_demux:src1_data -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:cp_data
	wire   [4:0] cmd_xbar_demux_src1_channel;                                                            // cmd_xbar_demux:src1_channel -> TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src2_endofpacket;                                                        // cmd_xbar_demux:src2_endofpacket -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                              // cmd_xbar_demux:src2_valid -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                      // cmd_xbar_demux:src2_startofpacket -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src2_data;                                                               // cmd_xbar_demux:src2_data -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:cp_data
	wire   [4:0] cmd_xbar_demux_src2_channel;                                                            // cmd_xbar_demux:src2_channel -> TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src3_endofpacket;                                                        // cmd_xbar_demux:src3_endofpacket -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                              // cmd_xbar_demux:src3_valid -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                      // cmd_xbar_demux:src3_startofpacket -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src3_data;                                                               // cmd_xbar_demux:src3_data -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:cp_data
	wire   [4:0] cmd_xbar_demux_src3_channel;                                                            // cmd_xbar_demux:src3_channel -> TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src4_endofpacket;                                                        // cmd_xbar_demux:src4_endofpacket -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                              // cmd_xbar_demux:src4_valid -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                      // cmd_xbar_demux:src4_startofpacket -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [86:0] cmd_xbar_demux_src4_data;                                                               // cmd_xbar_demux:src4_data -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [4:0] cmd_xbar_demux_src4_channel;                                                            // cmd_xbar_demux:src4_channel -> TEST_MEM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                        // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                              // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                      // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [86:0] rsp_xbar_demux_src0_data;                                                               // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [4:0] rsp_xbar_demux_src0_channel;                                                            // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                              // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                    // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                          // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                  // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [86:0] rsp_xbar_demux_001_src0_data;                                                           // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [4:0] rsp_xbar_demux_001_src0_channel;                                                        // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                          // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                    // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                          // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                  // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [86:0] rsp_xbar_demux_002_src0_data;                                                           // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [4:0] rsp_xbar_demux_002_src0_channel;                                                        // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                          // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                    // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                          // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                  // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [86:0] rsp_xbar_demux_003_src0_data;                                                           // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [4:0] rsp_xbar_demux_003_src0_channel;                                                        // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                          // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                    // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                          // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                  // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [86:0] rsp_xbar_demux_004_src0_data;                                                           // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [4:0] rsp_xbar_demux_004_src0_channel;                                                        // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                          // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                            // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                          // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [86:0] limiter_cmd_src_data;                                                                   // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [4:0] limiter_cmd_src_channel;                                                                // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                  // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                           // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                 // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                         // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [86:0] rsp_xbar_mux_src_data;                                                                  // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [4:0] rsp_xbar_mux_src_channel;                                                               // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                 // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         cmd_xbar_demux_src0_ready;                                                              // TEST_LED_TestReg_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire         id_router_src_endofpacket;                                                              // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                    // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                            // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [86:0] id_router_src_data;                                                                     // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [4:0] id_router_src_channel;                                                                  // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                    // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_demux_src1_ready;                                                              // TEST_REG0_TestReg_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire         id_router_001_src_endofpacket;                                                          // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                        // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [86:0] id_router_001_src_data;                                                                 // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [4:0] id_router_001_src_channel;                                                              // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_src2_ready;                                                              // TEST_REG1_TestReg_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	wire         id_router_002_src_endofpacket;                                                          // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                        // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [86:0] id_router_002_src_data;                                                                 // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [4:0] id_router_002_src_channel;                                                              // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_src3_ready;                                                              // TEST_REG2_TestReg_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src3_ready
	wire         id_router_003_src_endofpacket;                                                          // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                        // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [86:0] id_router_003_src_data;                                                                 // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [4:0] id_router_003_src_channel;                                                              // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_src4_ready;                                                              // TEST_MEM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src4_ready
	wire         id_router_004_src_endofpacket;                                                          // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                        // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [86:0] id_router_004_src_data;                                                                 // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [4:0] id_router_004_src_channel;                                                              // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire   [4:0] limiter_cmd_valid_data;                                                                 // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [9:0] sam9_host_events_irq;                                                                   // irq_synchronizer:sender_irq -> SAM9_HOST:inr_EVENTS_irq
	wire   [9:0] irq_synchronizer_receiver_irq;                                                          // irq_mapper:sender_irq -> irq_synchronizer:receiver_irq

	qsys_host_SAM9 sam9_host (
		.rso_MRST_reset       (sam9_host_mrst_reset),       //   MRST.reset
		.cso_MCLK_clk         (sam9_host_mclk_clk),         //   MCLK.clk
		.cso_H1CLK_clk        (),                           //  H1CLK.clk
		.cso_H2CLK_clk        (),                           //  H2CLK.clk
		.avm_M1_writedata     (sam9_host_m1_writedata),     //     M1.writedata
		.avm_M1_readdata      (sam9_host_m1_readdata),      //       .readdata
		.avm_M1_address       (sam9_host_m1_address),       //       .address
		.avm_M1_byteenable    (sam9_host_m1_byteenable),    //       .byteenable
		.avm_M1_write         (sam9_host_m1_write),         //       .write
		.avm_M1_read          (sam9_host_m1_read),          //       .read
		.avm_M1_begintransfer (sam9_host_m1_begintransfer), //       .begintransfer
		.avm_M1_readdatavalid (sam9_host_m1_readdatavalid), //       .readdatavalid
		.avm_M1_waitrequest   (sam9_host_m1_waitrequest),   //       .waitrequest
		.inr_EVENTS_irq       (sam9_host_events_irq),       // EVENTS.irq
		.coe_M1_RSTN          (m1_RSTN),                    // EXPORT.export
		.coe_M1_CLK           (m1_CLK),                     //       .export
		.coe_M1_ADDR          (m1_ADDR),                    //       .export
		.coe_M1_DATA          (m1_DATA),                    //       .export
		.coe_M1_CSN           (m1_CSN),                     //       .export
		.coe_M1_BEN           (m1_BEN),                     //       .export
		.coe_M1_RDN           (m1_RDN),                     //       .export
		.coe_M1_WRN           (m1_WRN),                     //       .export
		.coe_M1_WAITN         (m1_WAITN),                   //       .export
		.coe_M1_EINT          (m1_EINT)                     //       .export
	);

	qsys_test_LED test_led (
		.rsi_MRST_reset          (sam9_host_mrst_reset),                                        //    MRST.reset
		.csi_MCLK_clk            (sam9_host_mclk_clk),                                          //    MCLK.clk
		.avs_TestReg_readdata    (test_led_testreg_translator_avalon_anti_slave_0_readdata),    // TestReg.readdata
		.avs_TestReg_read        (test_led_testreg_translator_avalon_anti_slave_0_read),        //        .read
		.avs_TestReg_writedata   (test_led_testreg_translator_avalon_anti_slave_0_writedata),   //        .writedata
		.avs_TestReg_write       (test_led_testreg_translator_avalon_anti_slave_0_write),       //        .write
		.avs_TestReg_waitrequest (test_led_testreg_translator_avalon_anti_slave_0_waitrequest), //        .waitrequest
		.coe_LED_F0R             (led_F0R),                                                     //  EXPORT.export
		.coe_LED_F0G             (led_F0G),                                                     //        .export
		.coe_LED_F0B             (led_F0B),                                                     //        .export
		.coe_LED_F1R             (led_F1R),                                                     //        .export
		.coe_LED_F1G             (led_F1G),                                                     //        .export
		.coe_LED_F1B             (led_F1B),                                                     //        .export
		.coe_LED_F2R             (led_F2R),                                                     //        .export
		.coe_LED_F2G             (led_F2G),                                                     //        .export
		.coe_LED_F2B             (led_F2B),                                                     //        .export
		.coe_LED_F3R             (led_F3R),                                                     //        .export
		.coe_LED_F3G             (led_F3G),                                                     //        .export
		.coe_LED_F3B             (led_F3B)                                                      //        .export
	);

	qsys_test_RegRW test_reg0 (
		.csi_MCLK_clk            (sam9_host_mclk_clk),                                           //    MCLK.clk
		.rsi_MRST_reset          (sam9_host_mrst_reset),                                         //    MRST.reset
		.avs_TestReg_readdata    (test_reg0_testreg_translator_avalon_anti_slave_0_readdata),    // TestReg.readdata
		.avs_TestReg_read        (test_reg0_testreg_translator_avalon_anti_slave_0_read),        //        .read
		.avs_TestReg_writedata   (test_reg0_testreg_translator_avalon_anti_slave_0_writedata),   //        .writedata
		.avs_TestReg_write       (test_reg0_testreg_translator_avalon_anti_slave_0_write),       //        .write
		.avs_TestReg_waitrequest (test_reg0_testreg_translator_avalon_anti_slave_0_waitrequest)  //        .waitrequest
	);

	qsys_test_RegRW test_reg1 (
		.csi_MCLK_clk            (sam9_host_mclk_clk),                                           //    MCLK.clk
		.rsi_MRST_reset          (sam9_host_mrst_reset),                                         //    MRST.reset
		.avs_TestReg_readdata    (test_reg1_testreg_translator_avalon_anti_slave_0_readdata),    // TestReg.readdata
		.avs_TestReg_read        (test_reg1_testreg_translator_avalon_anti_slave_0_read),        //        .read
		.avs_TestReg_writedata   (test_reg1_testreg_translator_avalon_anti_slave_0_writedata),   //        .writedata
		.avs_TestReg_write       (test_reg1_testreg_translator_avalon_anti_slave_0_write),       //        .write
		.avs_TestReg_waitrequest (test_reg1_testreg_translator_avalon_anti_slave_0_waitrequest)  //        .waitrequest
	);

	qsys_test_RegRW test_reg2 (
		.csi_MCLK_clk            (sam9_host_mclk_clk),                                           //    MCLK.clk
		.rsi_MRST_reset          (sam9_host_mrst_reset),                                         //    MRST.reset
		.avs_TestReg_readdata    (test_reg2_testreg_translator_avalon_anti_slave_0_readdata),    // TestReg.readdata
		.avs_TestReg_read        (test_reg2_testreg_translator_avalon_anti_slave_0_read),        //        .read
		.avs_TestReg_writedata   (test_reg2_testreg_translator_avalon_anti_slave_0_writedata),   //        .writedata
		.avs_TestReg_write       (test_reg2_testreg_translator_avalon_anti_slave_0_write),       //        .write
		.avs_TestReg_waitrequest (test_reg2_testreg_translator_avalon_anti_slave_0_waitrequest)  //        .waitrequest
	);

	frontier_TEST_MEM test_mem (
		.clk        (sam9_host_mclk_clk),                                    //   clk1.clk
		.address    (test_mem_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (test_mem_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (test_mem_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (test_mem_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (test_mem_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (test_mem_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (test_mem_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (sam9_host_mrst_reset)                                   // reset1.reset
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (1),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sam9_host_m1_translator (
		.clk                   (sam9_host_mclk_clk),                                              //                       clk.clk
		.reset                 (sam9_host_mrst_reset),                                            //                     reset.reset
		.uav_address           (sam9_host_m1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (sam9_host_m1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (sam9_host_m1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (sam9_host_m1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (sam9_host_m1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (sam9_host_m1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (sam9_host_m1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (sam9_host_m1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (sam9_host_m1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (sam9_host_m1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (sam9_host_m1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (sam9_host_m1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (sam9_host_m1_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (sam9_host_m1_byteenable),                                         //                          .byteenable
		.av_begintransfer      (sam9_host_m1_begintransfer),                                      //                          .begintransfer
		.av_read               (sam9_host_m1_read),                                               //                          .read
		.av_readdata           (sam9_host_m1_readdata),                                           //                          .readdata
		.av_readdatavalid      (sam9_host_m1_readdatavalid),                                      //                          .readdatavalid
		.av_write              (sam9_host_m1_write),                                              //                          .write
		.av_writedata          (sam9_host_m1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                            //               (terminated)
		.av_chipselect         (1'b0),                                                            //               (terminated)
		.av_lock               (1'b0),                                                            //               (terminated)
		.av_debugaccess        (1'b0),                                                            //               (terminated)
		.uav_clken             (),                                                                //               (terminated)
		.av_clken              (1'b1)                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) test_led_testreg_translator (
		.clk                   (sam9_host_mclk_clk),                                                          //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                        //                    reset.reset
		.uav_address           (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (test_led_testreg_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (test_led_testreg_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (test_led_testreg_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (test_led_testreg_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (test_led_testreg_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_chipselect         (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) test_reg0_testreg_translator (
		.clk                   (sam9_host_mclk_clk),                                                           //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                         //                    reset.reset
		.uav_address           (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (test_reg0_testreg_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (test_reg0_testreg_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (test_reg0_testreg_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (test_reg0_testreg_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (test_reg0_testreg_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) test_reg1_testreg_translator (
		.clk                   (sam9_host_mclk_clk),                                                           //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                         //                    reset.reset
		.uav_address           (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (test_reg1_testreg_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (test_reg1_testreg_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (test_reg1_testreg_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (test_reg1_testreg_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (test_reg1_testreg_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) test_reg2_testreg_translator (
		.clk                   (sam9_host_mclk_clk),                                                           //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                         //                    reset.reset
		.uav_address           (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (test_reg2_testreg_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_read               (test_reg2_testreg_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (test_reg2_testreg_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (test_reg2_testreg_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (test_reg2_testreg_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_address            (),                                                                             //              (terminated)
		.av_begintransfer      (),                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) test_mem_s1_translator (
		.clk                   (sam9_host_mclk_clk),                                                     //                      clk.clk
		.reset                 (sam9_host_mrst_reset),                                                   //                    reset.reset
		.uav_address           (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (test_mem_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (test_mem_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (test_mem_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (test_mem_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (test_mem_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (test_mem_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (test_mem_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) test_reg2_testreg_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                                     //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                                   //       clk_reset.reset
		.m0_address              (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (test_reg2_testreg_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src3_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_src3_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_src3_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_src3_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src3_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src3_channel),                                                            //                .channel
		.rf_sink_ready           (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                                     //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                                   // clk_reset.reset
		.in_data           (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) test_mem_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                               //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                             //       clk_reset.reset
		.m0_address              (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (test_mem_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (test_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (test_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (test_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (test_mem_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (test_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src4_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_src4_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_src4_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_src4_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src4_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src4_channel),                                                      //                .channel
		.rf_sink_ready           (test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (test_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (test_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (test_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (test_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (test_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (test_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                               //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                             // clk_reset.reset
		.in_data           (test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (test_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (test_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) test_reg0_testreg_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                                     //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                                   //       clk_reset.reset
		.m0_address              (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (test_reg0_testreg_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                            //                .channel
		.rf_sink_ready           (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                                     //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                                   // clk_reset.reset
		.in_data           (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) test_reg1_testreg_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                                     //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                                   //       clk_reset.reset
		.m0_address              (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (test_reg1_testreg_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src2_ready),                                                              //              cp.ready
		.cp_valid                (cmd_xbar_demux_src2_valid),                                                              //                .valid
		.cp_data                 (cmd_xbar_demux_src2_data),                                                               //                .data
		.cp_startofpacket        (cmd_xbar_demux_src2_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src2_endofpacket),                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src2_channel),                                                            //                .channel
		.rf_sink_ready           (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                                     //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                                   // clk_reset.reset
		.in_data           (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) test_led_testreg_translator_avalon_universal_slave_0_agent (
		.clk                     (sam9_host_mclk_clk),                                                                    //             clk.clk
		.reset                   (sam9_host_mrst_reset),                                                                  //       clk_reset.reset
		.m0_address              (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (test_led_testreg_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (test_led_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (test_led_testreg_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (test_led_testreg_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (test_led_testreg_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (test_led_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                           //                .channel
		.rf_sink_ready           (test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (test_led_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (test_led_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (test_led_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (test_led_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (test_led_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (test_led_testreg_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sam9_host_mclk_clk),                                                                    //       clk.clk
		.reset             (sam9_host_mrst_reset),                                                                  // clk_reset.reset
		.in_data           (test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (test_led_testreg_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (test_led_testreg_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (86),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (78),
		.PKT_BURSTWRAP_L           (76),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (80),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7)
	) sam9_host_m1_translator_avalon_universal_master_0_agent (
		.clk              (sam9_host_mclk_clk),                                                       //       clk.clk
		.reset            (sam9_host_mrst_reset),                                                     // clk_reset.reset
		.av_address       (sam9_host_m1_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (sam9_host_m1_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (sam9_host_m1_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (sam9_host_m1_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (sam9_host_m1_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (sam9_host_m1_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (sam9_host_m1_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (sam9_host_m1_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (sam9_host_m1_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (sam9_host_m1_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (sam9_host_m1_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                    //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                     //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                  //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                     //          .ready
	);

	frontier_addr_router addr_router (
		.sink_ready         (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sam9_host_m1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                       //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_src_valid),                                                    //          .valid
		.src_data           (addr_router_src_data),                                                     //          .data
		.src_channel        (addr_router_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                               //          .endofpacket
	);

	frontier_id_router id_router (
		.sink_ready         (test_led_testreg_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (test_led_testreg_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (test_led_testreg_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (test_led_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (test_led_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                          //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                         //       src.ready
		.src_valid          (id_router_src_valid),                                                         //          .valid
		.src_data           (id_router_src_data),                                                          //          .data
		.src_channel        (id_router_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                    //          .endofpacket
	);

	frontier_id_router id_router_001 (
		.sink_ready         (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (test_reg0_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                           //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                      //       src.ready
		.src_valid          (id_router_001_src_valid),                                                      //          .valid
		.src_data           (id_router_001_src_data),                                                       //          .data
		.src_channel        (id_router_001_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router id_router_002 (
		.sink_ready         (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (test_reg1_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                           //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                      //       src.ready
		.src_valid          (id_router_002_src_valid),                                                      //          .valid
		.src_data           (id_router_002_src_data),                                                       //          .data
		.src_channel        (id_router_002_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router id_router_003 (
		.sink_ready         (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (test_reg2_testreg_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                           //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                      //       src.ready
		.src_valid          (id_router_003_src_valid),                                                      //          .valid
		.src_data           (id_router_003_src_data),                                                       //          .data
		.src_channel        (id_router_003_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                 //          .endofpacket
	);

	frontier_id_router id_router_004 (
		.sink_ready         (test_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (test_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (test_mem_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (test_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (test_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sam9_host_mclk_clk),                                                     //       clk.clk
		.reset              (sam9_host_mrst_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                //       src.ready
		.src_valid          (id_router_004_src_valid),                                                //          .valid
		.src_data           (id_router_004_src_data),                                                 //          .data
		.src_channel        (id_router_004_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                           //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (83),
		.PKT_TRANS_POSTED          (69),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (5),
		.VALID_WIDTH               (5),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (75),
		.PKT_BYTE_CNT_L            (73),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (sam9_host_mclk_clk),             //       clk.clk
		.reset                  (sam9_host_mrst_reset),           // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	frontier_cmd_xbar_demux cmd_xbar_demux (
		.clk                (sam9_host_mclk_clk),                //        clk.clk
		.reset              (sam9_host_mrst_reset),              //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket)    //           .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux (
		.clk                (sam9_host_mclk_clk),                //       clk.clk
		.reset              (sam9_host_mrst_reset),              // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (sam9_host_mclk_clk),                    //       clk.clk
		.reset              (sam9_host_mrst_reset),                  // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (sam9_host_mclk_clk),                    //       clk.clk
		.reset              (sam9_host_mrst_reset),                  // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (sam9_host_mclk_clk),                    //       clk.clk
		.reset              (sam9_host_mrst_reset),                  // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (sam9_host_mclk_clk),                    //       clk.clk
		.reset              (sam9_host_mrst_reset),                  // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	frontier_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (sam9_host_mclk_clk),                    //       clk.clk
		.reset               (sam9_host_mrst_reset),                  // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	frontier_irq_mapper irq_mapper (
		.clk        (sam9_host_mclk_clk),            //       clk.clk
		.reset      (sam9_host_mrst_reset),          // clk_reset.reset
		.sender_irq (irq_synchronizer_receiver_irq)  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (10)
	) irq_synchronizer (
		.receiver_clk   (sam9_host_mclk_clk),            //       receiver_clk.clk
		.sender_clk     (sam9_host_mclk_clk),            //         sender_clk.clk
		.receiver_reset (sam9_host_mrst_reset),          // receiver_clk_reset.reset
		.sender_reset   (sam9_host_mrst_reset),          //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq), //           receiver.irq
		.sender_irq     (sam9_host_events_irq)           //             sender.irq
	);

endmodule
